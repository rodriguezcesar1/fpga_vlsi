magic
tech scmos
timestamp 1608344865
<< ntransistor >>
rect 2701 4250 2703 4254
rect 2727 4246 2729 4250
rect 2732 4246 2734 4250
rect 2755 4242 2757 4246
rect 2887 4211 2889 4223
rect 2940 4211 2942 4223
rect 2727 4186 2729 4190
rect 2732 4186 2734 4190
rect 2679 4120 2681 4124
rect 2701 4120 2703 4124
rect 2727 4116 2729 4120
rect 2732 4116 2734 4120
rect 2755 4112 2757 4116
rect 2793 4081 2795 4093
rect 2846 4081 2848 4093
rect 2727 4056 2729 4060
rect 2732 4056 2734 4060
rect 1996 3715 1998 3719
rect 2001 3715 2003 3719
rect 2017 3715 2019 3719
rect 2033 3715 2035 3719
rect 2038 3715 2040 3719
rect 2059 3715 2061 3719
rect 2075 3715 2077 3719
rect 2091 3715 2093 3719
rect 2096 3715 2098 3719
rect 2112 3715 2114 3719
rect 2128 3715 2130 3719
rect 2133 3715 2135 3719
rect 2149 3715 2151 3719
rect 2165 3715 2167 3719
rect 2170 3715 2172 3719
rect 2191 3715 2193 3719
rect 2207 3715 2209 3719
rect 2223 3715 2225 3719
rect 2228 3715 2230 3719
rect 2244 3715 2246 3719
rect 2260 3715 2262 3719
rect 2265 3715 2267 3719
rect 2281 3715 2283 3719
rect 2297 3715 2299 3719
rect 2302 3715 2304 3719
rect 2323 3715 2325 3719
rect 2339 3715 2341 3719
rect 2355 3715 2357 3719
rect 2360 3715 2362 3719
rect 2376 3715 2378 3719
rect 2392 3715 2394 3719
rect 2397 3715 2399 3719
rect 2413 3715 2415 3719
rect 2429 3715 2431 3719
rect 2434 3715 2436 3719
rect 2455 3715 2457 3719
rect 2471 3715 2473 3719
rect 2487 3715 2489 3719
rect 2492 3715 2494 3719
rect 2508 3715 2510 3719
rect 2941 3715 2943 3719
rect 2946 3715 2948 3719
rect 2962 3715 2964 3719
rect 2978 3715 2980 3719
rect 2983 3715 2985 3719
rect 3004 3715 3006 3719
rect 3020 3715 3022 3719
rect 3036 3715 3038 3719
rect 3041 3715 3043 3719
rect 3057 3715 3059 3719
rect 3073 3715 3075 3719
rect 3078 3715 3080 3719
rect 3094 3715 3096 3719
rect 3110 3715 3112 3719
rect 3115 3715 3117 3719
rect 3136 3715 3138 3719
rect 3152 3715 3154 3719
rect 3168 3715 3170 3719
rect 3173 3715 3175 3719
rect 3189 3715 3191 3719
rect 3205 3715 3207 3719
rect 3210 3715 3212 3719
rect 3226 3715 3228 3719
rect 3242 3715 3244 3719
rect 3247 3715 3249 3719
rect 3268 3715 3270 3719
rect 3284 3715 3286 3719
rect 3300 3715 3302 3719
rect 3305 3715 3307 3719
rect 3321 3715 3323 3719
rect 3337 3715 3339 3719
rect 3342 3715 3344 3719
rect 3358 3715 3360 3719
rect 3374 3715 3376 3719
rect 3379 3715 3381 3719
rect 3400 3715 3402 3719
rect 3416 3715 3418 3719
rect 3432 3715 3434 3719
rect 3437 3715 3439 3719
rect 3453 3715 3455 3719
rect 1644 3682 1646 3686
rect 1649 3682 1651 3686
rect 1665 3682 1667 3686
rect 1681 3682 1683 3686
rect 1686 3682 1688 3686
rect 1707 3682 1709 3686
rect 1723 3682 1725 3686
rect 1739 3682 1741 3686
rect 1744 3682 1746 3686
rect 1760 3682 1762 3686
rect 2589 3682 2591 3686
rect 2594 3682 2596 3686
rect 2610 3682 2612 3686
rect 2626 3682 2628 3686
rect 2631 3682 2633 3686
rect 2652 3682 2654 3686
rect 2668 3682 2670 3686
rect 2684 3682 2686 3686
rect 2689 3682 2691 3686
rect 2705 3682 2707 3686
rect 1768 3645 1770 3649
rect 2175 3649 2177 3653
rect 2201 3645 2203 3649
rect 2206 3645 2208 3649
rect 2256 3649 2258 3653
rect 2282 3645 2284 3649
rect 2287 3645 2289 3649
rect 2229 3641 2231 3645
rect 1651 3636 1653 3640
rect 2001 3636 2003 3640
rect 2017 3636 2019 3640
rect 2033 3636 2035 3640
rect 2056 3636 2058 3640
rect 2061 3636 2063 3640
rect 2087 3636 2089 3640
rect 2108 3636 2110 3640
rect 2128 3636 2130 3640
rect 2133 3636 2135 3640
rect 2151 3636 2153 3640
rect 2310 3641 2312 3645
rect 2713 3645 2715 3649
rect 3120 3649 3122 3653
rect 3146 3645 3148 3649
rect 3151 3645 3153 3649
rect 3201 3649 3203 3653
rect 3227 3645 3229 3649
rect 3232 3645 3234 3649
rect 3174 3641 3176 3645
rect 2596 3636 2598 3640
rect 2946 3636 2948 3640
rect 2962 3636 2964 3640
rect 2978 3636 2980 3640
rect 3001 3636 3003 3640
rect 3006 3636 3008 3640
rect 3032 3636 3034 3640
rect 3053 3636 3055 3640
rect 3073 3636 3075 3640
rect 3078 3636 3080 3640
rect 3096 3636 3098 3640
rect 3255 3641 3257 3645
rect 2001 3590 2003 3594
rect 2017 3590 2019 3594
rect 2033 3590 2035 3594
rect 2056 3590 2058 3594
rect 2061 3590 2063 3594
rect 2087 3590 2089 3594
rect 2108 3590 2110 3594
rect 2128 3590 2130 3594
rect 2133 3590 2135 3594
rect 2151 3590 2153 3594
rect 1635 3580 1637 3584
rect 1651 3580 1653 3584
rect 1656 3580 1658 3584
rect 1672 3580 1674 3584
rect 1688 3580 1690 3584
rect 1709 3580 1711 3584
rect 1714 3580 1716 3584
rect 1730 3580 1732 3584
rect 1746 3580 1748 3584
rect 1751 3580 1753 3584
rect 2201 3589 2203 3593
rect 2206 3589 2208 3593
rect 2282 3589 2284 3593
rect 2287 3589 2289 3593
rect 2946 3590 2948 3594
rect 2962 3590 2964 3594
rect 2978 3590 2980 3594
rect 3001 3590 3003 3594
rect 3006 3590 3008 3594
rect 3032 3590 3034 3594
rect 3053 3590 3055 3594
rect 3073 3590 3075 3594
rect 3078 3590 3080 3594
rect 3096 3590 3098 3594
rect 2580 3580 2582 3584
rect 2596 3580 2598 3584
rect 2601 3580 2603 3584
rect 2617 3580 2619 3584
rect 2633 3580 2635 3584
rect 2654 3580 2656 3584
rect 2659 3580 2661 3584
rect 2675 3580 2677 3584
rect 2691 3580 2693 3584
rect 2696 3580 2698 3584
rect 3146 3589 3148 3593
rect 3151 3589 3153 3593
rect 3227 3589 3229 3593
rect 3232 3589 3234 3593
rect 2201 3513 2203 3517
rect 2206 3513 2208 3517
rect 2280 3517 2282 3521
rect 2306 3513 2308 3517
rect 2311 3513 2313 3517
rect 2229 3509 2231 3513
rect 2001 3504 2003 3508
rect 2017 3504 2019 3508
rect 2033 3504 2035 3508
rect 2056 3504 2058 3508
rect 2061 3504 2063 3508
rect 2087 3504 2089 3508
rect 2108 3504 2110 3508
rect 2128 3504 2130 3508
rect 2133 3504 2135 3508
rect 2151 3504 2153 3508
rect 2334 3509 2336 3513
rect 3146 3513 3148 3517
rect 3151 3513 3153 3517
rect 3225 3517 3227 3521
rect 3251 3513 3253 3517
rect 3256 3513 3258 3517
rect 3174 3509 3176 3513
rect 2946 3504 2948 3508
rect 2962 3504 2964 3508
rect 2978 3504 2980 3508
rect 3001 3504 3003 3508
rect 3006 3504 3008 3508
rect 3032 3504 3034 3508
rect 3053 3504 3055 3508
rect 3073 3504 3075 3508
rect 3078 3504 3080 3508
rect 3096 3504 3098 3508
rect 3279 3509 3281 3513
rect 2001 3458 2003 3462
rect 2017 3458 2019 3462
rect 2033 3458 2035 3462
rect 2056 3458 2058 3462
rect 2061 3458 2063 3462
rect 2087 3458 2089 3462
rect 2108 3458 2110 3462
rect 2128 3458 2130 3462
rect 2133 3458 2135 3462
rect 2151 3458 2153 3462
rect 2201 3458 2203 3462
rect 2206 3458 2208 3462
rect 2306 3458 2308 3462
rect 2311 3458 2313 3462
rect 2946 3458 2948 3462
rect 2962 3458 2964 3462
rect 2978 3458 2980 3462
rect 3001 3458 3003 3462
rect 3006 3458 3008 3462
rect 3032 3458 3034 3462
rect 3053 3458 3055 3462
rect 3073 3458 3075 3462
rect 3078 3458 3080 3462
rect 3096 3458 3098 3462
rect 3146 3458 3148 3462
rect 3151 3458 3153 3462
rect 3251 3458 3253 3462
rect 3256 3458 3258 3462
rect 2201 3381 2203 3385
rect 2206 3381 2208 3385
rect 2256 3385 2258 3389
rect 2282 3381 2284 3385
rect 2287 3381 2289 3385
rect 2346 3385 2348 3389
rect 2372 3381 2374 3385
rect 2377 3381 2379 3385
rect 2229 3377 2231 3381
rect 2001 3372 2003 3376
rect 2017 3372 2019 3376
rect 2033 3372 2035 3376
rect 2056 3372 2058 3376
rect 2061 3372 2063 3376
rect 2087 3372 2089 3376
rect 2108 3372 2110 3376
rect 2128 3372 2130 3376
rect 2133 3372 2135 3376
rect 2151 3372 2153 3376
rect 2310 3377 2312 3381
rect 2400 3377 2402 3381
rect 3146 3381 3148 3385
rect 3151 3381 3153 3385
rect 3201 3385 3203 3389
rect 3227 3381 3229 3385
rect 3232 3381 3234 3385
rect 3291 3385 3293 3389
rect 3317 3381 3319 3385
rect 3322 3381 3324 3385
rect 3174 3377 3176 3381
rect 2946 3372 2948 3376
rect 2962 3372 2964 3376
rect 2978 3372 2980 3376
rect 3001 3372 3003 3376
rect 3006 3372 3008 3376
rect 3032 3372 3034 3376
rect 3053 3372 3055 3376
rect 3073 3372 3075 3376
rect 3078 3372 3080 3376
rect 3096 3372 3098 3376
rect 3255 3377 3257 3381
rect 3345 3377 3347 3381
rect 2001 3326 2003 3330
rect 2017 3326 2019 3330
rect 2033 3326 2035 3330
rect 2056 3326 2058 3330
rect 2061 3326 2063 3330
rect 2087 3326 2089 3330
rect 2108 3326 2110 3330
rect 2128 3326 2130 3330
rect 2133 3326 2135 3330
rect 2151 3326 2153 3330
rect 2201 3323 2203 3327
rect 2206 3323 2208 3327
rect 2282 3323 2284 3327
rect 2287 3323 2289 3327
rect 2372 3323 2374 3327
rect 2377 3323 2379 3327
rect 2946 3326 2948 3330
rect 2962 3326 2964 3330
rect 2978 3326 2980 3330
rect 3001 3326 3003 3330
rect 3006 3326 3008 3330
rect 3032 3326 3034 3330
rect 3053 3326 3055 3330
rect 3073 3326 3075 3330
rect 3078 3326 3080 3330
rect 3096 3326 3098 3330
rect 3146 3323 3148 3327
rect 3151 3323 3153 3327
rect 3227 3323 3229 3327
rect 3232 3323 3234 3327
rect 3317 3323 3319 3327
rect 3322 3323 3324 3327
rect 2201 3249 2203 3253
rect 2206 3249 2208 3253
rect 2229 3245 2231 3249
rect 2001 3240 2003 3244
rect 2017 3240 2019 3244
rect 2033 3240 2035 3244
rect 2056 3240 2058 3244
rect 2061 3240 2063 3244
rect 2087 3240 2089 3244
rect 2108 3240 2110 3244
rect 2128 3240 2130 3244
rect 2133 3240 2135 3244
rect 2151 3240 2153 3244
rect 3146 3249 3148 3253
rect 3151 3249 3153 3253
rect 3174 3245 3176 3249
rect 2946 3240 2948 3244
rect 2962 3240 2964 3244
rect 2978 3240 2980 3244
rect 3001 3240 3003 3244
rect 3006 3240 3008 3244
rect 3032 3240 3034 3244
rect 3053 3240 3055 3244
rect 3073 3240 3075 3244
rect 3078 3240 3080 3244
rect 3096 3240 3098 3244
rect 2001 3194 2003 3198
rect 2017 3194 2019 3198
rect 2033 3194 2035 3198
rect 2056 3194 2058 3198
rect 2061 3194 2063 3198
rect 2087 3194 2089 3198
rect 2108 3194 2110 3198
rect 2128 3194 2130 3198
rect 2133 3194 2135 3198
rect 2151 3194 2153 3198
rect 2235 3194 2237 3198
rect 2253 3194 2255 3198
rect 2278 3194 2280 3198
rect 2294 3194 2296 3198
rect 2317 3194 2319 3198
rect 2322 3194 2324 3198
rect 2348 3194 2350 3198
rect 2369 3194 2371 3198
rect 2389 3194 2391 3198
rect 2394 3194 2396 3198
rect 2412 3194 2414 3198
rect 1512 3180 1514 3184
rect 1517 3180 1519 3184
rect 1533 3180 1535 3184
rect 1549 3180 1551 3184
rect 1554 3180 1556 3184
rect 1575 3180 1577 3184
rect 1591 3180 1593 3184
rect 1607 3180 1609 3184
rect 1612 3180 1614 3184
rect 1628 3180 1630 3184
rect 1644 3180 1646 3184
rect 1649 3180 1651 3184
rect 1665 3180 1667 3184
rect 1681 3180 1683 3184
rect 1686 3180 1688 3184
rect 1707 3180 1709 3184
rect 1723 3180 1725 3184
rect 1739 3180 1741 3184
rect 1744 3180 1746 3184
rect 1760 3180 1762 3184
rect 1776 3180 1778 3184
rect 1781 3180 1783 3184
rect 1797 3180 1799 3184
rect 1813 3180 1815 3184
rect 1818 3180 1820 3184
rect 1839 3180 1841 3184
rect 1855 3180 1857 3184
rect 1871 3180 1873 3184
rect 1876 3180 1878 3184
rect 1892 3180 1894 3184
rect 2201 3187 2203 3191
rect 2206 3187 2208 3191
rect 2946 3194 2948 3198
rect 2962 3194 2964 3198
rect 2978 3194 2980 3198
rect 3001 3194 3003 3198
rect 3006 3194 3008 3198
rect 3032 3194 3034 3198
rect 3053 3194 3055 3198
rect 3073 3194 3075 3198
rect 3078 3194 3080 3198
rect 3096 3194 3098 3198
rect 3180 3194 3182 3198
rect 3198 3194 3200 3198
rect 3223 3194 3225 3198
rect 3239 3194 3241 3198
rect 3262 3194 3264 3198
rect 3267 3194 3269 3198
rect 3293 3194 3295 3198
rect 3314 3194 3316 3198
rect 3334 3194 3336 3198
rect 3339 3194 3341 3198
rect 3357 3194 3359 3198
rect 2457 3180 2459 3184
rect 2462 3180 2464 3184
rect 2478 3180 2480 3184
rect 2494 3180 2496 3184
rect 2499 3180 2501 3184
rect 2520 3180 2522 3184
rect 2536 3180 2538 3184
rect 2552 3180 2554 3184
rect 2557 3180 2559 3184
rect 2573 3180 2575 3184
rect 2589 3180 2591 3184
rect 2594 3180 2596 3184
rect 2610 3180 2612 3184
rect 2626 3180 2628 3184
rect 2631 3180 2633 3184
rect 2652 3180 2654 3184
rect 2668 3180 2670 3184
rect 2684 3180 2686 3184
rect 2689 3180 2691 3184
rect 2705 3180 2707 3184
rect 2721 3180 2723 3184
rect 2726 3180 2728 3184
rect 2742 3180 2744 3184
rect 2758 3180 2760 3184
rect 2763 3180 2765 3184
rect 2784 3180 2786 3184
rect 2800 3180 2802 3184
rect 2816 3180 2818 3184
rect 2821 3180 2823 3184
rect 2837 3180 2839 3184
rect 3146 3187 3148 3191
rect 3151 3187 3153 3191
rect 1627 3136 1629 3140
rect 1651 3136 1653 3140
rect 2424 3138 2428 3140
rect 2572 3136 2574 3140
rect 2596 3136 2598 3140
rect 3369 3138 3373 3140
rect 1647 3123 1649 3127
rect 2592 3123 2594 3127
rect 1638 3109 1642 3111
rect 2583 3109 2587 3111
rect 1627 3100 1629 3104
rect 1651 3100 1653 3104
rect 2572 3100 2574 3104
rect 2596 3100 2598 3104
rect 2295 3068 2297 3072
rect 2300 3068 2302 3072
rect 2316 3068 2318 3072
rect 2332 3068 2334 3072
rect 2337 3068 2339 3072
rect 2358 3068 2360 3072
rect 2374 3068 2376 3072
rect 2390 3068 2392 3072
rect 2395 3068 2397 3072
rect 2411 3068 2413 3072
rect 3240 3068 3242 3072
rect 3245 3068 3247 3072
rect 3261 3068 3263 3072
rect 3277 3068 3279 3072
rect 3282 3068 3284 3072
rect 3303 3068 3305 3072
rect 3319 3068 3321 3072
rect 3335 3068 3337 3072
rect 3340 3068 3342 3072
rect 3356 3068 3358 3072
rect 1512 3038 1514 3042
rect 1517 3038 1519 3042
rect 1533 3038 1535 3042
rect 1549 3038 1551 3042
rect 1554 3038 1556 3042
rect 1575 3038 1577 3042
rect 1591 3038 1593 3042
rect 1607 3038 1609 3042
rect 1612 3038 1614 3042
rect 1628 3038 1630 3042
rect 1644 3038 1646 3042
rect 1649 3038 1651 3042
rect 1665 3038 1667 3042
rect 1681 3038 1683 3042
rect 1686 3038 1688 3042
rect 1707 3038 1709 3042
rect 1723 3038 1725 3042
rect 1739 3038 1741 3042
rect 1744 3038 1746 3042
rect 1760 3038 1762 3042
rect 1776 3038 1778 3042
rect 1781 3038 1783 3042
rect 1797 3038 1799 3042
rect 1813 3038 1815 3042
rect 1818 3038 1820 3042
rect 1839 3038 1841 3042
rect 1855 3038 1857 3042
rect 1871 3038 1873 3042
rect 1876 3038 1878 3042
rect 1892 3038 1894 3042
rect 2457 3038 2459 3042
rect 2462 3038 2464 3042
rect 2478 3038 2480 3042
rect 2494 3038 2496 3042
rect 2499 3038 2501 3042
rect 2520 3038 2522 3042
rect 2536 3038 2538 3042
rect 2552 3038 2554 3042
rect 2557 3038 2559 3042
rect 2573 3038 2575 3042
rect 2589 3038 2591 3042
rect 2594 3038 2596 3042
rect 2610 3038 2612 3042
rect 2626 3038 2628 3042
rect 2631 3038 2633 3042
rect 2652 3038 2654 3042
rect 2668 3038 2670 3042
rect 2684 3038 2686 3042
rect 2689 3038 2691 3042
rect 2705 3038 2707 3042
rect 2721 3038 2723 3042
rect 2726 3038 2728 3042
rect 2742 3038 2744 3042
rect 2758 3038 2760 3042
rect 2763 3038 2765 3042
rect 2784 3038 2786 3042
rect 2800 3038 2802 3042
rect 2816 3038 2818 3042
rect 2821 3038 2823 3042
rect 2837 3038 2839 3042
rect 2436 2992 2440 2994
rect 3381 2992 3385 2994
rect 2295 2982 2297 2986
rect 2300 2982 2302 2986
rect 2316 2982 2318 2986
rect 2332 2982 2334 2986
rect 2337 2982 2339 2986
rect 2358 2982 2360 2986
rect 2374 2982 2376 2986
rect 2390 2982 2392 2986
rect 2395 2982 2397 2986
rect 2411 2982 2413 2986
rect 3240 2982 3242 2986
rect 3245 2982 3247 2986
rect 3261 2982 3263 2986
rect 3277 2982 3279 2986
rect 3282 2982 3284 2986
rect 3303 2982 3305 2986
rect 3319 2982 3321 2986
rect 3335 2982 3337 2986
rect 3340 2982 3342 2986
rect 3356 2982 3358 2986
rect 1512 2952 1514 2956
rect 1517 2952 1519 2956
rect 1533 2952 1535 2956
rect 1549 2952 1551 2956
rect 1554 2952 1556 2956
rect 1575 2952 1577 2956
rect 1591 2952 1593 2956
rect 1607 2952 1609 2956
rect 1612 2952 1614 2956
rect 1628 2952 1630 2956
rect 1644 2952 1646 2956
rect 1649 2952 1651 2956
rect 1665 2952 1667 2956
rect 1681 2952 1683 2956
rect 1686 2952 1688 2956
rect 1707 2952 1709 2956
rect 1723 2952 1725 2956
rect 1739 2952 1741 2956
rect 1744 2952 1746 2956
rect 1760 2952 1762 2956
rect 1776 2952 1778 2956
rect 1781 2952 1783 2956
rect 1797 2952 1799 2956
rect 1813 2952 1815 2956
rect 1818 2952 1820 2956
rect 1839 2952 1841 2956
rect 1855 2952 1857 2956
rect 1871 2952 1873 2956
rect 1876 2952 1878 2956
rect 1892 2952 1894 2956
rect 2457 2952 2459 2956
rect 2462 2952 2464 2956
rect 2478 2952 2480 2956
rect 2494 2952 2496 2956
rect 2499 2952 2501 2956
rect 2520 2952 2522 2956
rect 2536 2952 2538 2956
rect 2552 2952 2554 2956
rect 2557 2952 2559 2956
rect 2573 2952 2575 2956
rect 2589 2952 2591 2956
rect 2594 2952 2596 2956
rect 2610 2952 2612 2956
rect 2626 2952 2628 2956
rect 2631 2952 2633 2956
rect 2652 2952 2654 2956
rect 2668 2952 2670 2956
rect 2684 2952 2686 2956
rect 2689 2952 2691 2956
rect 2705 2952 2707 2956
rect 2721 2952 2723 2956
rect 2726 2952 2728 2956
rect 2742 2952 2744 2956
rect 2758 2952 2760 2956
rect 2763 2952 2765 2956
rect 2784 2952 2786 2956
rect 2800 2952 2802 2956
rect 2816 2952 2818 2956
rect 2821 2952 2823 2956
rect 2837 2952 2839 2956
rect 1744 2908 1746 2912
rect 1768 2908 1770 2912
rect 2689 2908 2691 2912
rect 2713 2908 2715 2912
rect 1764 2897 1766 2901
rect 2709 2897 2711 2901
rect 1755 2883 1759 2885
rect 2700 2883 2704 2885
rect 1744 2874 1746 2878
rect 1768 2874 1770 2878
rect 2689 2874 2691 2878
rect 2713 2874 2715 2878
rect 1512 2812 1514 2816
rect 1517 2812 1519 2816
rect 1533 2812 1535 2816
rect 1549 2812 1551 2816
rect 1554 2812 1556 2816
rect 1575 2812 1577 2816
rect 1591 2812 1593 2816
rect 1607 2812 1609 2816
rect 1612 2812 1614 2816
rect 1628 2812 1630 2816
rect 1644 2812 1646 2816
rect 1649 2812 1651 2816
rect 1665 2812 1667 2816
rect 1681 2812 1683 2816
rect 1686 2812 1688 2816
rect 1707 2812 1709 2816
rect 1723 2812 1725 2816
rect 1739 2812 1741 2816
rect 1744 2812 1746 2816
rect 1760 2812 1762 2816
rect 1776 2812 1778 2816
rect 1781 2812 1783 2816
rect 1797 2812 1799 2816
rect 1813 2812 1815 2816
rect 1818 2812 1820 2816
rect 1839 2812 1841 2816
rect 1855 2812 1857 2816
rect 1871 2812 1873 2816
rect 1876 2812 1878 2816
rect 1892 2812 1894 2816
rect 2457 2812 2459 2816
rect 2462 2812 2464 2816
rect 2478 2812 2480 2816
rect 2494 2812 2496 2816
rect 2499 2812 2501 2816
rect 2520 2812 2522 2816
rect 2536 2812 2538 2816
rect 2552 2812 2554 2816
rect 2557 2812 2559 2816
rect 2573 2812 2575 2816
rect 2589 2812 2591 2816
rect 2594 2812 2596 2816
rect 2610 2812 2612 2816
rect 2626 2812 2628 2816
rect 2631 2812 2633 2816
rect 2652 2812 2654 2816
rect 2668 2812 2670 2816
rect 2684 2812 2686 2816
rect 2689 2812 2691 2816
rect 2705 2812 2707 2816
rect 2721 2812 2723 2816
rect 2726 2812 2728 2816
rect 2742 2812 2744 2816
rect 2758 2812 2760 2816
rect 2763 2812 2765 2816
rect 2784 2812 2786 2816
rect 2800 2812 2802 2816
rect 2816 2812 2818 2816
rect 2821 2812 2823 2816
rect 2837 2812 2839 2816
rect 1996 2733 1998 2737
rect 2001 2733 2003 2737
rect 2017 2733 2019 2737
rect 2033 2733 2035 2737
rect 2038 2733 2040 2737
rect 2059 2733 2061 2737
rect 2075 2733 2077 2737
rect 2091 2733 2093 2737
rect 2096 2733 2098 2737
rect 2112 2733 2114 2737
rect 2128 2733 2130 2737
rect 2133 2733 2135 2737
rect 2149 2733 2151 2737
rect 2165 2733 2167 2737
rect 2170 2733 2172 2737
rect 2191 2733 2193 2737
rect 2207 2733 2209 2737
rect 2223 2733 2225 2737
rect 2228 2733 2230 2737
rect 2244 2733 2246 2737
rect 2260 2733 2262 2737
rect 2265 2733 2267 2737
rect 2281 2733 2283 2737
rect 2297 2733 2299 2737
rect 2302 2733 2304 2737
rect 2323 2733 2325 2737
rect 2339 2733 2341 2737
rect 2355 2733 2357 2737
rect 2360 2733 2362 2737
rect 2376 2733 2378 2737
rect 2392 2733 2394 2737
rect 2397 2733 2399 2737
rect 2413 2733 2415 2737
rect 2429 2733 2431 2737
rect 2434 2733 2436 2737
rect 2455 2733 2457 2737
rect 2471 2733 2473 2737
rect 2487 2733 2489 2737
rect 2492 2733 2494 2737
rect 2508 2733 2510 2737
rect 2941 2733 2943 2737
rect 2946 2733 2948 2737
rect 2962 2733 2964 2737
rect 2978 2733 2980 2737
rect 2983 2733 2985 2737
rect 3004 2733 3006 2737
rect 3020 2733 3022 2737
rect 3036 2733 3038 2737
rect 3041 2733 3043 2737
rect 3057 2733 3059 2737
rect 3073 2733 3075 2737
rect 3078 2733 3080 2737
rect 3094 2733 3096 2737
rect 3110 2733 3112 2737
rect 3115 2733 3117 2737
rect 3136 2733 3138 2737
rect 3152 2733 3154 2737
rect 3168 2733 3170 2737
rect 3173 2733 3175 2737
rect 3189 2733 3191 2737
rect 3205 2733 3207 2737
rect 3210 2733 3212 2737
rect 3226 2733 3228 2737
rect 3242 2733 3244 2737
rect 3247 2733 3249 2737
rect 3268 2733 3270 2737
rect 3284 2733 3286 2737
rect 3300 2733 3302 2737
rect 3305 2733 3307 2737
rect 3321 2733 3323 2737
rect 3337 2733 3339 2737
rect 3342 2733 3344 2737
rect 3358 2733 3360 2737
rect 3374 2733 3376 2737
rect 3379 2733 3381 2737
rect 3400 2733 3402 2737
rect 3416 2733 3418 2737
rect 3432 2733 3434 2737
rect 3437 2733 3439 2737
rect 3453 2733 3455 2737
rect 1644 2700 1646 2704
rect 1649 2700 1651 2704
rect 1665 2700 1667 2704
rect 1681 2700 1683 2704
rect 1686 2700 1688 2704
rect 1707 2700 1709 2704
rect 1723 2700 1725 2704
rect 1739 2700 1741 2704
rect 1744 2700 1746 2704
rect 1760 2700 1762 2704
rect 2589 2700 2591 2704
rect 2594 2700 2596 2704
rect 2610 2700 2612 2704
rect 2626 2700 2628 2704
rect 2631 2700 2633 2704
rect 2652 2700 2654 2704
rect 2668 2700 2670 2704
rect 2684 2700 2686 2704
rect 2689 2700 2691 2704
rect 2705 2700 2707 2704
rect 1768 2663 1770 2667
rect 2175 2667 2177 2671
rect 2201 2663 2203 2667
rect 2206 2663 2208 2667
rect 2256 2667 2258 2671
rect 2282 2663 2284 2667
rect 2287 2663 2289 2667
rect 2229 2659 2231 2663
rect 1651 2654 1653 2658
rect 2001 2654 2003 2658
rect 2017 2654 2019 2658
rect 2033 2654 2035 2658
rect 2056 2654 2058 2658
rect 2061 2654 2063 2658
rect 2087 2654 2089 2658
rect 2108 2654 2110 2658
rect 2128 2654 2130 2658
rect 2133 2654 2135 2658
rect 2151 2654 2153 2658
rect 2310 2659 2312 2663
rect 2713 2663 2715 2667
rect 3120 2667 3122 2671
rect 3146 2663 3148 2667
rect 3151 2663 3153 2667
rect 3201 2667 3203 2671
rect 3227 2663 3229 2667
rect 3232 2663 3234 2667
rect 3174 2659 3176 2663
rect 2596 2654 2598 2658
rect 2946 2654 2948 2658
rect 2962 2654 2964 2658
rect 2978 2654 2980 2658
rect 3001 2654 3003 2658
rect 3006 2654 3008 2658
rect 3032 2654 3034 2658
rect 3053 2654 3055 2658
rect 3073 2654 3075 2658
rect 3078 2654 3080 2658
rect 3096 2654 3098 2658
rect 3255 2659 3257 2663
rect 2001 2608 2003 2612
rect 2017 2608 2019 2612
rect 2033 2608 2035 2612
rect 2056 2608 2058 2612
rect 2061 2608 2063 2612
rect 2087 2608 2089 2612
rect 2108 2608 2110 2612
rect 2128 2608 2130 2612
rect 2133 2608 2135 2612
rect 2151 2608 2153 2612
rect 1635 2598 1637 2602
rect 1651 2598 1653 2602
rect 1656 2598 1658 2602
rect 1672 2598 1674 2602
rect 1688 2598 1690 2602
rect 1709 2598 1711 2602
rect 1714 2598 1716 2602
rect 1730 2598 1732 2602
rect 1746 2598 1748 2602
rect 1751 2598 1753 2602
rect 2201 2607 2203 2611
rect 2206 2607 2208 2611
rect 2282 2607 2284 2611
rect 2287 2607 2289 2611
rect 2946 2608 2948 2612
rect 2962 2608 2964 2612
rect 2978 2608 2980 2612
rect 3001 2608 3003 2612
rect 3006 2608 3008 2612
rect 3032 2608 3034 2612
rect 3053 2608 3055 2612
rect 3073 2608 3075 2612
rect 3078 2608 3080 2612
rect 3096 2608 3098 2612
rect 2580 2598 2582 2602
rect 2596 2598 2598 2602
rect 2601 2598 2603 2602
rect 2617 2598 2619 2602
rect 2633 2598 2635 2602
rect 2654 2598 2656 2602
rect 2659 2598 2661 2602
rect 2675 2598 2677 2602
rect 2691 2598 2693 2602
rect 2696 2598 2698 2602
rect 3146 2607 3148 2611
rect 3151 2607 3153 2611
rect 3227 2607 3229 2611
rect 3232 2607 3234 2611
rect 2201 2531 2203 2535
rect 2206 2531 2208 2535
rect 2280 2535 2282 2539
rect 2306 2531 2308 2535
rect 2311 2531 2313 2535
rect 2229 2527 2231 2531
rect 2001 2522 2003 2526
rect 2017 2522 2019 2526
rect 2033 2522 2035 2526
rect 2056 2522 2058 2526
rect 2061 2522 2063 2526
rect 2087 2522 2089 2526
rect 2108 2522 2110 2526
rect 2128 2522 2130 2526
rect 2133 2522 2135 2526
rect 2151 2522 2153 2526
rect 2334 2527 2336 2531
rect 3146 2531 3148 2535
rect 3151 2531 3153 2535
rect 3225 2535 3227 2539
rect 3251 2531 3253 2535
rect 3256 2531 3258 2535
rect 3174 2527 3176 2531
rect 2946 2522 2948 2526
rect 2962 2522 2964 2526
rect 2978 2522 2980 2526
rect 3001 2522 3003 2526
rect 3006 2522 3008 2526
rect 3032 2522 3034 2526
rect 3053 2522 3055 2526
rect 3073 2522 3075 2526
rect 3078 2522 3080 2526
rect 3096 2522 3098 2526
rect 3279 2527 3281 2531
rect 2001 2476 2003 2480
rect 2017 2476 2019 2480
rect 2033 2476 2035 2480
rect 2056 2476 2058 2480
rect 2061 2476 2063 2480
rect 2087 2476 2089 2480
rect 2108 2476 2110 2480
rect 2128 2476 2130 2480
rect 2133 2476 2135 2480
rect 2151 2476 2153 2480
rect 2201 2476 2203 2480
rect 2206 2476 2208 2480
rect 2306 2476 2308 2480
rect 2311 2476 2313 2480
rect 2946 2476 2948 2480
rect 2962 2476 2964 2480
rect 2978 2476 2980 2480
rect 3001 2476 3003 2480
rect 3006 2476 3008 2480
rect 3032 2476 3034 2480
rect 3053 2476 3055 2480
rect 3073 2476 3075 2480
rect 3078 2476 3080 2480
rect 3096 2476 3098 2480
rect 3146 2476 3148 2480
rect 3151 2476 3153 2480
rect 3251 2476 3253 2480
rect 3256 2476 3258 2480
rect 2201 2399 2203 2403
rect 2206 2399 2208 2403
rect 2256 2403 2258 2407
rect 2282 2399 2284 2403
rect 2287 2399 2289 2403
rect 2346 2403 2348 2407
rect 2372 2399 2374 2403
rect 2377 2399 2379 2403
rect 2229 2395 2231 2399
rect 2001 2390 2003 2394
rect 2017 2390 2019 2394
rect 2033 2390 2035 2394
rect 2056 2390 2058 2394
rect 2061 2390 2063 2394
rect 2087 2390 2089 2394
rect 2108 2390 2110 2394
rect 2128 2390 2130 2394
rect 2133 2390 2135 2394
rect 2151 2390 2153 2394
rect 2310 2395 2312 2399
rect 2400 2395 2402 2399
rect 3146 2399 3148 2403
rect 3151 2399 3153 2403
rect 3201 2403 3203 2407
rect 3227 2399 3229 2403
rect 3232 2399 3234 2403
rect 3291 2403 3293 2407
rect 3317 2399 3319 2403
rect 3322 2399 3324 2403
rect 3174 2395 3176 2399
rect 2946 2390 2948 2394
rect 2962 2390 2964 2394
rect 2978 2390 2980 2394
rect 3001 2390 3003 2394
rect 3006 2390 3008 2394
rect 3032 2390 3034 2394
rect 3053 2390 3055 2394
rect 3073 2390 3075 2394
rect 3078 2390 3080 2394
rect 3096 2390 3098 2394
rect 3255 2395 3257 2399
rect 3345 2395 3347 2399
rect 2001 2344 2003 2348
rect 2017 2344 2019 2348
rect 2033 2344 2035 2348
rect 2056 2344 2058 2348
rect 2061 2344 2063 2348
rect 2087 2344 2089 2348
rect 2108 2344 2110 2348
rect 2128 2344 2130 2348
rect 2133 2344 2135 2348
rect 2151 2344 2153 2348
rect 2201 2341 2203 2345
rect 2206 2341 2208 2345
rect 2282 2341 2284 2345
rect 2287 2341 2289 2345
rect 2372 2341 2374 2345
rect 2377 2341 2379 2345
rect 2946 2344 2948 2348
rect 2962 2344 2964 2348
rect 2978 2344 2980 2348
rect 3001 2344 3003 2348
rect 3006 2344 3008 2348
rect 3032 2344 3034 2348
rect 3053 2344 3055 2348
rect 3073 2344 3075 2348
rect 3078 2344 3080 2348
rect 3096 2344 3098 2348
rect 3146 2341 3148 2345
rect 3151 2341 3153 2345
rect 3227 2341 3229 2345
rect 3232 2341 3234 2345
rect 3317 2341 3319 2345
rect 3322 2341 3324 2345
rect 2201 2267 2203 2271
rect 2206 2267 2208 2271
rect 2229 2263 2231 2267
rect 2001 2258 2003 2262
rect 2017 2258 2019 2262
rect 2033 2258 2035 2262
rect 2056 2258 2058 2262
rect 2061 2258 2063 2262
rect 2087 2258 2089 2262
rect 2108 2258 2110 2262
rect 2128 2258 2130 2262
rect 2133 2258 2135 2262
rect 2151 2258 2153 2262
rect 3146 2267 3148 2271
rect 3151 2267 3153 2271
rect 3174 2263 3176 2267
rect 2946 2258 2948 2262
rect 2962 2258 2964 2262
rect 2978 2258 2980 2262
rect 3001 2258 3003 2262
rect 3006 2258 3008 2262
rect 3032 2258 3034 2262
rect 3053 2258 3055 2262
rect 3073 2258 3075 2262
rect 3078 2258 3080 2262
rect 3096 2258 3098 2262
rect 2001 2212 2003 2216
rect 2017 2212 2019 2216
rect 2033 2212 2035 2216
rect 2056 2212 2058 2216
rect 2061 2212 2063 2216
rect 2087 2212 2089 2216
rect 2108 2212 2110 2216
rect 2128 2212 2130 2216
rect 2133 2212 2135 2216
rect 2151 2212 2153 2216
rect 2235 2212 2237 2216
rect 2253 2212 2255 2216
rect 2278 2212 2280 2216
rect 2294 2212 2296 2216
rect 2317 2212 2319 2216
rect 2322 2212 2324 2216
rect 2348 2212 2350 2216
rect 2369 2212 2371 2216
rect 2389 2212 2391 2216
rect 2394 2212 2396 2216
rect 2412 2212 2414 2216
rect 1512 2198 1514 2202
rect 1517 2198 1519 2202
rect 1533 2198 1535 2202
rect 1549 2198 1551 2202
rect 1554 2198 1556 2202
rect 1575 2198 1577 2202
rect 1591 2198 1593 2202
rect 1607 2198 1609 2202
rect 1612 2198 1614 2202
rect 1628 2198 1630 2202
rect 1644 2198 1646 2202
rect 1649 2198 1651 2202
rect 1665 2198 1667 2202
rect 1681 2198 1683 2202
rect 1686 2198 1688 2202
rect 1707 2198 1709 2202
rect 1723 2198 1725 2202
rect 1739 2198 1741 2202
rect 1744 2198 1746 2202
rect 1760 2198 1762 2202
rect 1776 2198 1778 2202
rect 1781 2198 1783 2202
rect 1797 2198 1799 2202
rect 1813 2198 1815 2202
rect 1818 2198 1820 2202
rect 1839 2198 1841 2202
rect 1855 2198 1857 2202
rect 1871 2198 1873 2202
rect 1876 2198 1878 2202
rect 1892 2198 1894 2202
rect 2201 2205 2203 2209
rect 2206 2205 2208 2209
rect 2946 2212 2948 2216
rect 2962 2212 2964 2216
rect 2978 2212 2980 2216
rect 3001 2212 3003 2216
rect 3006 2212 3008 2216
rect 3032 2212 3034 2216
rect 3053 2212 3055 2216
rect 3073 2212 3075 2216
rect 3078 2212 3080 2216
rect 3096 2212 3098 2216
rect 3180 2212 3182 2216
rect 3198 2212 3200 2216
rect 3223 2212 3225 2216
rect 3239 2212 3241 2216
rect 3262 2212 3264 2216
rect 3267 2212 3269 2216
rect 3293 2212 3295 2216
rect 3314 2212 3316 2216
rect 3334 2212 3336 2216
rect 3339 2212 3341 2216
rect 3357 2212 3359 2216
rect 2457 2198 2459 2202
rect 2462 2198 2464 2202
rect 2478 2198 2480 2202
rect 2494 2198 2496 2202
rect 2499 2198 2501 2202
rect 2520 2198 2522 2202
rect 2536 2198 2538 2202
rect 2552 2198 2554 2202
rect 2557 2198 2559 2202
rect 2573 2198 2575 2202
rect 2589 2198 2591 2202
rect 2594 2198 2596 2202
rect 2610 2198 2612 2202
rect 2626 2198 2628 2202
rect 2631 2198 2633 2202
rect 2652 2198 2654 2202
rect 2668 2198 2670 2202
rect 2684 2198 2686 2202
rect 2689 2198 2691 2202
rect 2705 2198 2707 2202
rect 2721 2198 2723 2202
rect 2726 2198 2728 2202
rect 2742 2198 2744 2202
rect 2758 2198 2760 2202
rect 2763 2198 2765 2202
rect 2784 2198 2786 2202
rect 2800 2198 2802 2202
rect 2816 2198 2818 2202
rect 2821 2198 2823 2202
rect 2837 2198 2839 2202
rect 3146 2205 3148 2209
rect 3151 2205 3153 2209
rect 1627 2154 1629 2158
rect 1651 2154 1653 2158
rect 2424 2156 2428 2158
rect 2572 2154 2574 2158
rect 2596 2154 2598 2158
rect 3369 2156 3373 2158
rect 1647 2141 1649 2145
rect 2592 2141 2594 2145
rect 1638 2127 1642 2129
rect 2583 2127 2587 2129
rect 1627 2118 1629 2122
rect 1651 2118 1653 2122
rect 2572 2118 2574 2122
rect 2596 2118 2598 2122
rect 2295 2086 2297 2090
rect 2300 2086 2302 2090
rect 2316 2086 2318 2090
rect 2332 2086 2334 2090
rect 2337 2086 2339 2090
rect 2358 2086 2360 2090
rect 2374 2086 2376 2090
rect 2390 2086 2392 2090
rect 2395 2086 2397 2090
rect 2411 2086 2413 2090
rect 3240 2086 3242 2090
rect 3245 2086 3247 2090
rect 3261 2086 3263 2090
rect 3277 2086 3279 2090
rect 3282 2086 3284 2090
rect 3303 2086 3305 2090
rect 3319 2086 3321 2090
rect 3335 2086 3337 2090
rect 3340 2086 3342 2090
rect 3356 2086 3358 2090
rect 1512 2056 1514 2060
rect 1517 2056 1519 2060
rect 1533 2056 1535 2060
rect 1549 2056 1551 2060
rect 1554 2056 1556 2060
rect 1575 2056 1577 2060
rect 1591 2056 1593 2060
rect 1607 2056 1609 2060
rect 1612 2056 1614 2060
rect 1628 2056 1630 2060
rect 1644 2056 1646 2060
rect 1649 2056 1651 2060
rect 1665 2056 1667 2060
rect 1681 2056 1683 2060
rect 1686 2056 1688 2060
rect 1707 2056 1709 2060
rect 1723 2056 1725 2060
rect 1739 2056 1741 2060
rect 1744 2056 1746 2060
rect 1760 2056 1762 2060
rect 1776 2056 1778 2060
rect 1781 2056 1783 2060
rect 1797 2056 1799 2060
rect 1813 2056 1815 2060
rect 1818 2056 1820 2060
rect 1839 2056 1841 2060
rect 1855 2056 1857 2060
rect 1871 2056 1873 2060
rect 1876 2056 1878 2060
rect 1892 2056 1894 2060
rect 2457 2056 2459 2060
rect 2462 2056 2464 2060
rect 2478 2056 2480 2060
rect 2494 2056 2496 2060
rect 2499 2056 2501 2060
rect 2520 2056 2522 2060
rect 2536 2056 2538 2060
rect 2552 2056 2554 2060
rect 2557 2056 2559 2060
rect 2573 2056 2575 2060
rect 2589 2056 2591 2060
rect 2594 2056 2596 2060
rect 2610 2056 2612 2060
rect 2626 2056 2628 2060
rect 2631 2056 2633 2060
rect 2652 2056 2654 2060
rect 2668 2056 2670 2060
rect 2684 2056 2686 2060
rect 2689 2056 2691 2060
rect 2705 2056 2707 2060
rect 2721 2056 2723 2060
rect 2726 2056 2728 2060
rect 2742 2056 2744 2060
rect 2758 2056 2760 2060
rect 2763 2056 2765 2060
rect 2784 2056 2786 2060
rect 2800 2056 2802 2060
rect 2816 2056 2818 2060
rect 2821 2056 2823 2060
rect 2837 2056 2839 2060
rect 2436 2010 2440 2012
rect 3381 2010 3385 2012
rect 2295 2000 2297 2004
rect 2300 2000 2302 2004
rect 2316 2000 2318 2004
rect 2332 2000 2334 2004
rect 2337 2000 2339 2004
rect 2358 2000 2360 2004
rect 2374 2000 2376 2004
rect 2390 2000 2392 2004
rect 2395 2000 2397 2004
rect 2411 2000 2413 2004
rect 3240 2000 3242 2004
rect 3245 2000 3247 2004
rect 3261 2000 3263 2004
rect 3277 2000 3279 2004
rect 3282 2000 3284 2004
rect 3303 2000 3305 2004
rect 3319 2000 3321 2004
rect 3335 2000 3337 2004
rect 3340 2000 3342 2004
rect 3356 2000 3358 2004
rect 1512 1970 1514 1974
rect 1517 1970 1519 1974
rect 1533 1970 1535 1974
rect 1549 1970 1551 1974
rect 1554 1970 1556 1974
rect 1575 1970 1577 1974
rect 1591 1970 1593 1974
rect 1607 1970 1609 1974
rect 1612 1970 1614 1974
rect 1628 1970 1630 1974
rect 1644 1970 1646 1974
rect 1649 1970 1651 1974
rect 1665 1970 1667 1974
rect 1681 1970 1683 1974
rect 1686 1970 1688 1974
rect 1707 1970 1709 1974
rect 1723 1970 1725 1974
rect 1739 1970 1741 1974
rect 1744 1970 1746 1974
rect 1760 1970 1762 1974
rect 1776 1970 1778 1974
rect 1781 1970 1783 1974
rect 1797 1970 1799 1974
rect 1813 1970 1815 1974
rect 1818 1970 1820 1974
rect 1839 1970 1841 1974
rect 1855 1970 1857 1974
rect 1871 1970 1873 1974
rect 1876 1970 1878 1974
rect 1892 1970 1894 1974
rect 2457 1970 2459 1974
rect 2462 1970 2464 1974
rect 2478 1970 2480 1974
rect 2494 1970 2496 1974
rect 2499 1970 2501 1974
rect 2520 1970 2522 1974
rect 2536 1970 2538 1974
rect 2552 1970 2554 1974
rect 2557 1970 2559 1974
rect 2573 1970 2575 1974
rect 2589 1970 2591 1974
rect 2594 1970 2596 1974
rect 2610 1970 2612 1974
rect 2626 1970 2628 1974
rect 2631 1970 2633 1974
rect 2652 1970 2654 1974
rect 2668 1970 2670 1974
rect 2684 1970 2686 1974
rect 2689 1970 2691 1974
rect 2705 1970 2707 1974
rect 2721 1970 2723 1974
rect 2726 1970 2728 1974
rect 2742 1970 2744 1974
rect 2758 1970 2760 1974
rect 2763 1970 2765 1974
rect 2784 1970 2786 1974
rect 2800 1970 2802 1974
rect 2816 1970 2818 1974
rect 2821 1970 2823 1974
rect 2837 1970 2839 1974
rect 1744 1926 1746 1930
rect 1768 1926 1770 1930
rect 2689 1926 2691 1930
rect 2713 1926 2715 1930
rect 1764 1915 1766 1919
rect 2709 1915 2711 1919
rect 1755 1901 1759 1903
rect 2700 1901 2704 1903
rect 1744 1892 1746 1896
rect 1768 1892 1770 1896
rect 2689 1892 2691 1896
rect 2713 1892 2715 1896
rect 1512 1830 1514 1834
rect 1517 1830 1519 1834
rect 1533 1830 1535 1834
rect 1549 1830 1551 1834
rect 1554 1830 1556 1834
rect 1575 1830 1577 1834
rect 1591 1830 1593 1834
rect 1607 1830 1609 1834
rect 1612 1830 1614 1834
rect 1628 1830 1630 1834
rect 1644 1830 1646 1834
rect 1649 1830 1651 1834
rect 1665 1830 1667 1834
rect 1681 1830 1683 1834
rect 1686 1830 1688 1834
rect 1707 1830 1709 1834
rect 1723 1830 1725 1834
rect 1739 1830 1741 1834
rect 1744 1830 1746 1834
rect 1760 1830 1762 1834
rect 1776 1830 1778 1834
rect 1781 1830 1783 1834
rect 1797 1830 1799 1834
rect 1813 1830 1815 1834
rect 1818 1830 1820 1834
rect 1839 1830 1841 1834
rect 1855 1830 1857 1834
rect 1871 1830 1873 1834
rect 1876 1830 1878 1834
rect 1892 1830 1894 1834
rect 2457 1830 2459 1834
rect 2462 1830 2464 1834
rect 2478 1830 2480 1834
rect 2494 1830 2496 1834
rect 2499 1830 2501 1834
rect 2520 1830 2522 1834
rect 2536 1830 2538 1834
rect 2552 1830 2554 1834
rect 2557 1830 2559 1834
rect 2573 1830 2575 1834
rect 2589 1830 2591 1834
rect 2594 1830 2596 1834
rect 2610 1830 2612 1834
rect 2626 1830 2628 1834
rect 2631 1830 2633 1834
rect 2652 1830 2654 1834
rect 2668 1830 2670 1834
rect 2684 1830 2686 1834
rect 2689 1830 2691 1834
rect 2705 1830 2707 1834
rect 2721 1830 2723 1834
rect 2726 1830 2728 1834
rect 2742 1830 2744 1834
rect 2758 1830 2760 1834
rect 2763 1830 2765 1834
rect 2784 1830 2786 1834
rect 2800 1830 2802 1834
rect 2816 1830 2818 1834
rect 2821 1830 2823 1834
rect 2837 1830 2839 1834
<< ptransistor >>
rect 2701 4268 2703 4276
rect 2727 4262 2729 4270
rect 2732 4262 2734 4270
rect 2755 4268 2757 4276
rect 2887 4243 2889 4273
rect 2940 4243 2942 4273
rect 2727 4166 2729 4174
rect 2732 4166 2734 4174
rect 2679 4138 2681 4146
rect 2701 4138 2703 4146
rect 2727 4132 2729 4140
rect 2732 4132 2734 4140
rect 2755 4138 2757 4146
rect 2793 4113 2795 4143
rect 2846 4113 2848 4143
rect 2727 4036 2729 4044
rect 2732 4036 2734 4044
rect 1996 3738 1998 3746
rect 2001 3738 2003 3746
rect 2017 3738 2019 3746
rect 2033 3738 2035 3746
rect 2038 3738 2040 3746
rect 2059 3738 2061 3746
rect 2075 3738 2077 3746
rect 2091 3738 2093 3746
rect 2096 3738 2098 3746
rect 2112 3738 2114 3746
rect 2128 3738 2130 3746
rect 2133 3738 2135 3746
rect 2149 3738 2151 3746
rect 2165 3738 2167 3746
rect 2170 3738 2172 3746
rect 2191 3738 2193 3746
rect 2207 3738 2209 3746
rect 2223 3738 2225 3746
rect 2228 3738 2230 3746
rect 2244 3738 2246 3746
rect 2260 3738 2262 3746
rect 2265 3738 2267 3746
rect 2281 3738 2283 3746
rect 2297 3738 2299 3746
rect 2302 3738 2304 3746
rect 2323 3738 2325 3746
rect 2339 3738 2341 3746
rect 2355 3738 2357 3746
rect 2360 3738 2362 3746
rect 2376 3738 2378 3746
rect 2392 3738 2394 3746
rect 2397 3738 2399 3746
rect 2413 3738 2415 3746
rect 2429 3738 2431 3746
rect 2434 3738 2436 3746
rect 2455 3738 2457 3746
rect 2471 3738 2473 3746
rect 2487 3738 2489 3746
rect 2492 3738 2494 3746
rect 2508 3738 2510 3746
rect 2941 3738 2943 3746
rect 2946 3738 2948 3746
rect 2962 3738 2964 3746
rect 2978 3738 2980 3746
rect 2983 3738 2985 3746
rect 3004 3738 3006 3746
rect 3020 3738 3022 3746
rect 3036 3738 3038 3746
rect 3041 3738 3043 3746
rect 3057 3738 3059 3746
rect 3073 3738 3075 3746
rect 3078 3738 3080 3746
rect 3094 3738 3096 3746
rect 3110 3738 3112 3746
rect 3115 3738 3117 3746
rect 3136 3738 3138 3746
rect 3152 3738 3154 3746
rect 3168 3738 3170 3746
rect 3173 3738 3175 3746
rect 3189 3738 3191 3746
rect 3205 3738 3207 3746
rect 3210 3738 3212 3746
rect 3226 3738 3228 3746
rect 3242 3738 3244 3746
rect 3247 3738 3249 3746
rect 3268 3738 3270 3746
rect 3284 3738 3286 3746
rect 3300 3738 3302 3746
rect 3305 3738 3307 3746
rect 3321 3738 3323 3746
rect 3337 3738 3339 3746
rect 3342 3738 3344 3746
rect 3358 3738 3360 3746
rect 3374 3738 3376 3746
rect 3379 3738 3381 3746
rect 3400 3738 3402 3746
rect 3416 3738 3418 3746
rect 3432 3738 3434 3746
rect 3437 3738 3439 3746
rect 3453 3738 3455 3746
rect 1644 3705 1646 3713
rect 1649 3705 1651 3713
rect 1665 3705 1667 3713
rect 1681 3705 1683 3713
rect 1686 3705 1688 3713
rect 1707 3705 1709 3713
rect 1723 3705 1725 3713
rect 1739 3705 1741 3713
rect 1744 3705 1746 3713
rect 1760 3705 1762 3713
rect 2589 3705 2591 3713
rect 2594 3705 2596 3713
rect 2610 3705 2612 3713
rect 2626 3705 2628 3713
rect 2631 3705 2633 3713
rect 2652 3705 2654 3713
rect 2668 3705 2670 3713
rect 2684 3705 2686 3713
rect 2689 3705 2691 3713
rect 2705 3705 2707 3713
rect 2175 3667 2177 3675
rect 2001 3654 2003 3662
rect 2017 3654 2019 3662
rect 2033 3654 2035 3662
rect 2056 3654 2058 3662
rect 2061 3654 2063 3662
rect 2087 3654 2089 3662
rect 2108 3654 2110 3662
rect 2128 3654 2130 3662
rect 2133 3654 2135 3662
rect 2151 3654 2153 3662
rect 2201 3661 2203 3669
rect 2206 3661 2208 3669
rect 2229 3667 2231 3675
rect 2256 3667 2258 3675
rect 2282 3661 2284 3669
rect 2287 3661 2289 3669
rect 2310 3667 2312 3675
rect 3120 3667 3122 3675
rect 2946 3654 2948 3662
rect 2962 3654 2964 3662
rect 2978 3654 2980 3662
rect 3001 3654 3003 3662
rect 3006 3654 3008 3662
rect 3032 3654 3034 3662
rect 3053 3654 3055 3662
rect 3073 3654 3075 3662
rect 3078 3654 3080 3662
rect 3096 3654 3098 3662
rect 3146 3661 3148 3669
rect 3151 3661 3153 3669
rect 3174 3667 3176 3675
rect 3201 3667 3203 3675
rect 3227 3661 3229 3669
rect 3232 3661 3234 3669
rect 3255 3667 3257 3675
rect 1635 3603 1637 3611
rect 1651 3603 1653 3611
rect 1656 3603 1658 3611
rect 1672 3603 1674 3611
rect 1688 3603 1690 3611
rect 1709 3603 1711 3611
rect 1714 3603 1716 3611
rect 1730 3603 1732 3611
rect 1746 3603 1748 3611
rect 1751 3603 1753 3611
rect 2580 3603 2582 3611
rect 2596 3603 2598 3611
rect 2601 3603 2603 3611
rect 2617 3603 2619 3611
rect 2633 3603 2635 3611
rect 2654 3603 2656 3611
rect 2659 3603 2661 3611
rect 2675 3603 2677 3611
rect 2691 3603 2693 3611
rect 2696 3603 2698 3611
rect 2001 3568 2003 3576
rect 2017 3568 2019 3576
rect 2033 3568 2035 3576
rect 2056 3568 2058 3576
rect 2061 3568 2063 3576
rect 2087 3568 2089 3576
rect 2108 3568 2110 3576
rect 2128 3568 2130 3576
rect 2133 3568 2135 3576
rect 2151 3568 2153 3576
rect 2201 3569 2203 3577
rect 2206 3569 2208 3577
rect 2282 3569 2284 3577
rect 2287 3569 2289 3577
rect 2946 3568 2948 3576
rect 2962 3568 2964 3576
rect 2978 3568 2980 3576
rect 3001 3568 3003 3576
rect 3006 3568 3008 3576
rect 3032 3568 3034 3576
rect 3053 3568 3055 3576
rect 3073 3568 3075 3576
rect 3078 3568 3080 3576
rect 3096 3568 3098 3576
rect 3146 3569 3148 3577
rect 3151 3569 3153 3577
rect 3227 3569 3229 3577
rect 3232 3569 3234 3577
rect 2001 3522 2003 3530
rect 2017 3522 2019 3530
rect 2033 3522 2035 3530
rect 2056 3522 2058 3530
rect 2061 3522 2063 3530
rect 2087 3522 2089 3530
rect 2108 3522 2110 3530
rect 2128 3522 2130 3530
rect 2133 3522 2135 3530
rect 2151 3522 2153 3530
rect 2201 3529 2203 3537
rect 2206 3529 2208 3537
rect 2229 3535 2231 3543
rect 2280 3535 2282 3543
rect 2306 3529 2308 3537
rect 2311 3529 2313 3537
rect 2334 3535 2336 3543
rect 2946 3522 2948 3530
rect 2962 3522 2964 3530
rect 2978 3522 2980 3530
rect 3001 3522 3003 3530
rect 3006 3522 3008 3530
rect 3032 3522 3034 3530
rect 3053 3522 3055 3530
rect 3073 3522 3075 3530
rect 3078 3522 3080 3530
rect 3096 3522 3098 3530
rect 3146 3529 3148 3537
rect 3151 3529 3153 3537
rect 3174 3535 3176 3543
rect 3225 3535 3227 3543
rect 3251 3529 3253 3537
rect 3256 3529 3258 3537
rect 3279 3535 3281 3543
rect 2001 3436 2003 3444
rect 2017 3436 2019 3444
rect 2033 3436 2035 3444
rect 2056 3436 2058 3444
rect 2061 3436 2063 3444
rect 2087 3436 2089 3444
rect 2108 3436 2110 3444
rect 2128 3436 2130 3444
rect 2133 3436 2135 3444
rect 2151 3436 2153 3444
rect 2201 3438 2203 3446
rect 2206 3438 2208 3446
rect 2306 3438 2308 3446
rect 2311 3438 2313 3446
rect 2946 3436 2948 3444
rect 2962 3436 2964 3444
rect 2978 3436 2980 3444
rect 3001 3436 3003 3444
rect 3006 3436 3008 3444
rect 3032 3436 3034 3444
rect 3053 3436 3055 3444
rect 3073 3436 3075 3444
rect 3078 3436 3080 3444
rect 3096 3436 3098 3444
rect 3146 3438 3148 3446
rect 3151 3438 3153 3446
rect 3251 3438 3253 3446
rect 3256 3438 3258 3446
rect 2001 3390 2003 3398
rect 2017 3390 2019 3398
rect 2033 3390 2035 3398
rect 2056 3390 2058 3398
rect 2061 3390 2063 3398
rect 2087 3390 2089 3398
rect 2108 3390 2110 3398
rect 2128 3390 2130 3398
rect 2133 3390 2135 3398
rect 2151 3390 2153 3398
rect 2201 3397 2203 3405
rect 2206 3397 2208 3405
rect 2229 3403 2231 3411
rect 2256 3403 2258 3411
rect 2282 3397 2284 3405
rect 2287 3397 2289 3405
rect 2310 3403 2312 3411
rect 2346 3403 2348 3411
rect 2372 3397 2374 3405
rect 2377 3397 2379 3405
rect 2400 3403 2402 3411
rect 2946 3390 2948 3398
rect 2962 3390 2964 3398
rect 2978 3390 2980 3398
rect 3001 3390 3003 3398
rect 3006 3390 3008 3398
rect 3032 3390 3034 3398
rect 3053 3390 3055 3398
rect 3073 3390 3075 3398
rect 3078 3390 3080 3398
rect 3096 3390 3098 3398
rect 3146 3397 3148 3405
rect 3151 3397 3153 3405
rect 3174 3403 3176 3411
rect 3201 3403 3203 3411
rect 3227 3397 3229 3405
rect 3232 3397 3234 3405
rect 3255 3403 3257 3411
rect 3291 3403 3293 3411
rect 3317 3397 3319 3405
rect 3322 3397 3324 3405
rect 3345 3403 3347 3411
rect 2001 3304 2003 3312
rect 2017 3304 2019 3312
rect 2033 3304 2035 3312
rect 2056 3304 2058 3312
rect 2061 3304 2063 3312
rect 2087 3304 2089 3312
rect 2108 3304 2110 3312
rect 2128 3304 2130 3312
rect 2133 3304 2135 3312
rect 2151 3304 2153 3312
rect 2201 3303 2203 3311
rect 2206 3303 2208 3311
rect 2282 3303 2284 3311
rect 2287 3303 2289 3311
rect 2372 3303 2374 3311
rect 2377 3303 2379 3311
rect 2946 3304 2948 3312
rect 2962 3304 2964 3312
rect 2978 3304 2980 3312
rect 3001 3304 3003 3312
rect 3006 3304 3008 3312
rect 3032 3304 3034 3312
rect 3053 3304 3055 3312
rect 3073 3304 3075 3312
rect 3078 3304 3080 3312
rect 3096 3304 3098 3312
rect 3146 3303 3148 3311
rect 3151 3303 3153 3311
rect 3227 3303 3229 3311
rect 3232 3303 3234 3311
rect 3317 3303 3319 3311
rect 3322 3303 3324 3311
rect 2001 3258 2003 3266
rect 2017 3258 2019 3266
rect 2033 3258 2035 3266
rect 2056 3258 2058 3266
rect 2061 3258 2063 3266
rect 2087 3258 2089 3266
rect 2108 3258 2110 3266
rect 2128 3258 2130 3266
rect 2133 3258 2135 3266
rect 2151 3258 2153 3266
rect 2201 3265 2203 3273
rect 2206 3265 2208 3273
rect 2229 3271 2231 3279
rect 2946 3258 2948 3266
rect 2962 3258 2964 3266
rect 2978 3258 2980 3266
rect 3001 3258 3003 3266
rect 3006 3258 3008 3266
rect 3032 3258 3034 3266
rect 3053 3258 3055 3266
rect 3073 3258 3075 3266
rect 3078 3258 3080 3266
rect 3096 3258 3098 3266
rect 3146 3265 3148 3273
rect 3151 3265 3153 3273
rect 3174 3271 3176 3279
rect 1512 3203 1514 3211
rect 1517 3203 1519 3211
rect 1533 3203 1535 3211
rect 1549 3203 1551 3211
rect 1554 3203 1556 3211
rect 1575 3203 1577 3211
rect 1591 3203 1593 3211
rect 1607 3203 1609 3211
rect 1612 3203 1614 3211
rect 1628 3203 1630 3211
rect 1644 3203 1646 3211
rect 1649 3203 1651 3211
rect 1665 3203 1667 3211
rect 1681 3203 1683 3211
rect 1686 3203 1688 3211
rect 1707 3203 1709 3211
rect 1723 3203 1725 3211
rect 1739 3203 1741 3211
rect 1744 3203 1746 3211
rect 1760 3203 1762 3211
rect 1776 3203 1778 3211
rect 1781 3203 1783 3211
rect 1797 3203 1799 3211
rect 1813 3203 1815 3211
rect 1818 3203 1820 3211
rect 1839 3203 1841 3211
rect 1855 3203 1857 3211
rect 1871 3203 1873 3211
rect 1876 3203 1878 3211
rect 1892 3203 1894 3211
rect 2457 3203 2459 3211
rect 2462 3203 2464 3211
rect 2478 3203 2480 3211
rect 2494 3203 2496 3211
rect 2499 3203 2501 3211
rect 2520 3203 2522 3211
rect 2536 3203 2538 3211
rect 2552 3203 2554 3211
rect 2557 3203 2559 3211
rect 2573 3203 2575 3211
rect 2589 3203 2591 3211
rect 2594 3203 2596 3211
rect 2610 3203 2612 3211
rect 2626 3203 2628 3211
rect 2631 3203 2633 3211
rect 2652 3203 2654 3211
rect 2668 3203 2670 3211
rect 2684 3203 2686 3211
rect 2689 3203 2691 3211
rect 2705 3203 2707 3211
rect 2721 3203 2723 3211
rect 2726 3203 2728 3211
rect 2742 3203 2744 3211
rect 2758 3203 2760 3211
rect 2763 3203 2765 3211
rect 2784 3203 2786 3211
rect 2800 3203 2802 3211
rect 2816 3203 2818 3211
rect 2821 3203 2823 3211
rect 2837 3203 2839 3211
rect 2001 3172 2003 3180
rect 2017 3172 2019 3180
rect 2033 3172 2035 3180
rect 2056 3172 2058 3180
rect 2061 3172 2063 3180
rect 2087 3172 2089 3180
rect 2108 3172 2110 3180
rect 2128 3172 2130 3180
rect 2133 3172 2135 3180
rect 2151 3172 2153 3180
rect 2201 3167 2203 3175
rect 2206 3167 2208 3175
rect 2235 3172 2237 3180
rect 2253 3172 2255 3180
rect 2278 3172 2280 3180
rect 2294 3172 2296 3180
rect 2317 3172 2319 3180
rect 2322 3172 2324 3180
rect 2348 3172 2350 3180
rect 2369 3172 2371 3180
rect 2389 3172 2391 3180
rect 2394 3172 2396 3180
rect 2412 3172 2414 3180
rect 2946 3172 2948 3180
rect 2962 3172 2964 3180
rect 2978 3172 2980 3180
rect 3001 3172 3003 3180
rect 3006 3172 3008 3180
rect 3032 3172 3034 3180
rect 3053 3172 3055 3180
rect 3073 3172 3075 3180
rect 3078 3172 3080 3180
rect 3096 3172 3098 3180
rect 3146 3167 3148 3175
rect 3151 3167 3153 3175
rect 3180 3172 3182 3180
rect 3198 3172 3200 3180
rect 3223 3172 3225 3180
rect 3239 3172 3241 3180
rect 3262 3172 3264 3180
rect 3267 3172 3269 3180
rect 3293 3172 3295 3180
rect 3314 3172 3316 3180
rect 3334 3172 3336 3180
rect 3339 3172 3341 3180
rect 3357 3172 3359 3180
rect 2295 3091 2297 3099
rect 2300 3091 2302 3099
rect 2316 3091 2318 3099
rect 2332 3091 2334 3099
rect 2337 3091 2339 3099
rect 2358 3091 2360 3099
rect 2374 3091 2376 3099
rect 2390 3091 2392 3099
rect 2395 3091 2397 3099
rect 2411 3091 2413 3099
rect 3240 3091 3242 3099
rect 3245 3091 3247 3099
rect 3261 3091 3263 3099
rect 3277 3091 3279 3099
rect 3282 3091 3284 3099
rect 3303 3091 3305 3099
rect 3319 3091 3321 3099
rect 3335 3091 3337 3099
rect 3340 3091 3342 3099
rect 3356 3091 3358 3099
rect 1512 3061 1514 3069
rect 1517 3061 1519 3069
rect 1533 3061 1535 3069
rect 1549 3061 1551 3069
rect 1554 3061 1556 3069
rect 1575 3061 1577 3069
rect 1591 3061 1593 3069
rect 1607 3061 1609 3069
rect 1612 3061 1614 3069
rect 1628 3061 1630 3069
rect 1644 3061 1646 3069
rect 1649 3061 1651 3069
rect 1665 3061 1667 3069
rect 1681 3061 1683 3069
rect 1686 3061 1688 3069
rect 1707 3061 1709 3069
rect 1723 3061 1725 3069
rect 1739 3061 1741 3069
rect 1744 3061 1746 3069
rect 1760 3061 1762 3069
rect 1776 3061 1778 3069
rect 1781 3061 1783 3069
rect 1797 3061 1799 3069
rect 1813 3061 1815 3069
rect 1818 3061 1820 3069
rect 1839 3061 1841 3069
rect 1855 3061 1857 3069
rect 1871 3061 1873 3069
rect 1876 3061 1878 3069
rect 1892 3061 1894 3069
rect 2457 3061 2459 3069
rect 2462 3061 2464 3069
rect 2478 3061 2480 3069
rect 2494 3061 2496 3069
rect 2499 3061 2501 3069
rect 2520 3061 2522 3069
rect 2536 3061 2538 3069
rect 2552 3061 2554 3069
rect 2557 3061 2559 3069
rect 2573 3061 2575 3069
rect 2589 3061 2591 3069
rect 2594 3061 2596 3069
rect 2610 3061 2612 3069
rect 2626 3061 2628 3069
rect 2631 3061 2633 3069
rect 2652 3061 2654 3069
rect 2668 3061 2670 3069
rect 2684 3061 2686 3069
rect 2689 3061 2691 3069
rect 2705 3061 2707 3069
rect 2721 3061 2723 3069
rect 2726 3061 2728 3069
rect 2742 3061 2744 3069
rect 2758 3061 2760 3069
rect 2763 3061 2765 3069
rect 2784 3061 2786 3069
rect 2800 3061 2802 3069
rect 2816 3061 2818 3069
rect 2821 3061 2823 3069
rect 2837 3061 2839 3069
rect 2295 3005 2297 3013
rect 2300 3005 2302 3013
rect 2316 3005 2318 3013
rect 2332 3005 2334 3013
rect 2337 3005 2339 3013
rect 2358 3005 2360 3013
rect 2374 3005 2376 3013
rect 2390 3005 2392 3013
rect 2395 3005 2397 3013
rect 2411 3005 2413 3013
rect 3240 3005 3242 3013
rect 3245 3005 3247 3013
rect 3261 3005 3263 3013
rect 3277 3005 3279 3013
rect 3282 3005 3284 3013
rect 3303 3005 3305 3013
rect 3319 3005 3321 3013
rect 3335 3005 3337 3013
rect 3340 3005 3342 3013
rect 3356 3005 3358 3013
rect 1512 2975 1514 2983
rect 1517 2975 1519 2983
rect 1533 2975 1535 2983
rect 1549 2975 1551 2983
rect 1554 2975 1556 2983
rect 1575 2975 1577 2983
rect 1591 2975 1593 2983
rect 1607 2975 1609 2983
rect 1612 2975 1614 2983
rect 1628 2975 1630 2983
rect 1644 2975 1646 2983
rect 1649 2975 1651 2983
rect 1665 2975 1667 2983
rect 1681 2975 1683 2983
rect 1686 2975 1688 2983
rect 1707 2975 1709 2983
rect 1723 2975 1725 2983
rect 1739 2975 1741 2983
rect 1744 2975 1746 2983
rect 1760 2975 1762 2983
rect 1776 2975 1778 2983
rect 1781 2975 1783 2983
rect 1797 2975 1799 2983
rect 1813 2975 1815 2983
rect 1818 2975 1820 2983
rect 1839 2975 1841 2983
rect 1855 2975 1857 2983
rect 1871 2975 1873 2983
rect 1876 2975 1878 2983
rect 1892 2975 1894 2983
rect 2457 2975 2459 2983
rect 2462 2975 2464 2983
rect 2478 2975 2480 2983
rect 2494 2975 2496 2983
rect 2499 2975 2501 2983
rect 2520 2975 2522 2983
rect 2536 2975 2538 2983
rect 2552 2975 2554 2983
rect 2557 2975 2559 2983
rect 2573 2975 2575 2983
rect 2589 2975 2591 2983
rect 2594 2975 2596 2983
rect 2610 2975 2612 2983
rect 2626 2975 2628 2983
rect 2631 2975 2633 2983
rect 2652 2975 2654 2983
rect 2668 2975 2670 2983
rect 2684 2975 2686 2983
rect 2689 2975 2691 2983
rect 2705 2975 2707 2983
rect 2721 2975 2723 2983
rect 2726 2975 2728 2983
rect 2742 2975 2744 2983
rect 2758 2975 2760 2983
rect 2763 2975 2765 2983
rect 2784 2975 2786 2983
rect 2800 2975 2802 2983
rect 2816 2975 2818 2983
rect 2821 2975 2823 2983
rect 2837 2975 2839 2983
rect 1512 2835 1514 2843
rect 1517 2835 1519 2843
rect 1533 2835 1535 2843
rect 1549 2835 1551 2843
rect 1554 2835 1556 2843
rect 1575 2835 1577 2843
rect 1591 2835 1593 2843
rect 1607 2835 1609 2843
rect 1612 2835 1614 2843
rect 1628 2835 1630 2843
rect 1644 2835 1646 2843
rect 1649 2835 1651 2843
rect 1665 2835 1667 2843
rect 1681 2835 1683 2843
rect 1686 2835 1688 2843
rect 1707 2835 1709 2843
rect 1723 2835 1725 2843
rect 1739 2835 1741 2843
rect 1744 2835 1746 2843
rect 1760 2835 1762 2843
rect 1776 2835 1778 2843
rect 1781 2835 1783 2843
rect 1797 2835 1799 2843
rect 1813 2835 1815 2843
rect 1818 2835 1820 2843
rect 1839 2835 1841 2843
rect 1855 2835 1857 2843
rect 1871 2835 1873 2843
rect 1876 2835 1878 2843
rect 1892 2835 1894 2843
rect 2457 2835 2459 2843
rect 2462 2835 2464 2843
rect 2478 2835 2480 2843
rect 2494 2835 2496 2843
rect 2499 2835 2501 2843
rect 2520 2835 2522 2843
rect 2536 2835 2538 2843
rect 2552 2835 2554 2843
rect 2557 2835 2559 2843
rect 2573 2835 2575 2843
rect 2589 2835 2591 2843
rect 2594 2835 2596 2843
rect 2610 2835 2612 2843
rect 2626 2835 2628 2843
rect 2631 2835 2633 2843
rect 2652 2835 2654 2843
rect 2668 2835 2670 2843
rect 2684 2835 2686 2843
rect 2689 2835 2691 2843
rect 2705 2835 2707 2843
rect 2721 2835 2723 2843
rect 2726 2835 2728 2843
rect 2742 2835 2744 2843
rect 2758 2835 2760 2843
rect 2763 2835 2765 2843
rect 2784 2835 2786 2843
rect 2800 2835 2802 2843
rect 2816 2835 2818 2843
rect 2821 2835 2823 2843
rect 2837 2835 2839 2843
rect 1996 2756 1998 2764
rect 2001 2756 2003 2764
rect 2017 2756 2019 2764
rect 2033 2756 2035 2764
rect 2038 2756 2040 2764
rect 2059 2756 2061 2764
rect 2075 2756 2077 2764
rect 2091 2756 2093 2764
rect 2096 2756 2098 2764
rect 2112 2756 2114 2764
rect 2128 2756 2130 2764
rect 2133 2756 2135 2764
rect 2149 2756 2151 2764
rect 2165 2756 2167 2764
rect 2170 2756 2172 2764
rect 2191 2756 2193 2764
rect 2207 2756 2209 2764
rect 2223 2756 2225 2764
rect 2228 2756 2230 2764
rect 2244 2756 2246 2764
rect 2260 2756 2262 2764
rect 2265 2756 2267 2764
rect 2281 2756 2283 2764
rect 2297 2756 2299 2764
rect 2302 2756 2304 2764
rect 2323 2756 2325 2764
rect 2339 2756 2341 2764
rect 2355 2756 2357 2764
rect 2360 2756 2362 2764
rect 2376 2756 2378 2764
rect 2392 2756 2394 2764
rect 2397 2756 2399 2764
rect 2413 2756 2415 2764
rect 2429 2756 2431 2764
rect 2434 2756 2436 2764
rect 2455 2756 2457 2764
rect 2471 2756 2473 2764
rect 2487 2756 2489 2764
rect 2492 2756 2494 2764
rect 2508 2756 2510 2764
rect 2941 2756 2943 2764
rect 2946 2756 2948 2764
rect 2962 2756 2964 2764
rect 2978 2756 2980 2764
rect 2983 2756 2985 2764
rect 3004 2756 3006 2764
rect 3020 2756 3022 2764
rect 3036 2756 3038 2764
rect 3041 2756 3043 2764
rect 3057 2756 3059 2764
rect 3073 2756 3075 2764
rect 3078 2756 3080 2764
rect 3094 2756 3096 2764
rect 3110 2756 3112 2764
rect 3115 2756 3117 2764
rect 3136 2756 3138 2764
rect 3152 2756 3154 2764
rect 3168 2756 3170 2764
rect 3173 2756 3175 2764
rect 3189 2756 3191 2764
rect 3205 2756 3207 2764
rect 3210 2756 3212 2764
rect 3226 2756 3228 2764
rect 3242 2756 3244 2764
rect 3247 2756 3249 2764
rect 3268 2756 3270 2764
rect 3284 2756 3286 2764
rect 3300 2756 3302 2764
rect 3305 2756 3307 2764
rect 3321 2756 3323 2764
rect 3337 2756 3339 2764
rect 3342 2756 3344 2764
rect 3358 2756 3360 2764
rect 3374 2756 3376 2764
rect 3379 2756 3381 2764
rect 3400 2756 3402 2764
rect 3416 2756 3418 2764
rect 3432 2756 3434 2764
rect 3437 2756 3439 2764
rect 3453 2756 3455 2764
rect 1644 2723 1646 2731
rect 1649 2723 1651 2731
rect 1665 2723 1667 2731
rect 1681 2723 1683 2731
rect 1686 2723 1688 2731
rect 1707 2723 1709 2731
rect 1723 2723 1725 2731
rect 1739 2723 1741 2731
rect 1744 2723 1746 2731
rect 1760 2723 1762 2731
rect 2589 2723 2591 2731
rect 2594 2723 2596 2731
rect 2610 2723 2612 2731
rect 2626 2723 2628 2731
rect 2631 2723 2633 2731
rect 2652 2723 2654 2731
rect 2668 2723 2670 2731
rect 2684 2723 2686 2731
rect 2689 2723 2691 2731
rect 2705 2723 2707 2731
rect 2175 2685 2177 2693
rect 2001 2672 2003 2680
rect 2017 2672 2019 2680
rect 2033 2672 2035 2680
rect 2056 2672 2058 2680
rect 2061 2672 2063 2680
rect 2087 2672 2089 2680
rect 2108 2672 2110 2680
rect 2128 2672 2130 2680
rect 2133 2672 2135 2680
rect 2151 2672 2153 2680
rect 2201 2679 2203 2687
rect 2206 2679 2208 2687
rect 2229 2685 2231 2693
rect 2256 2685 2258 2693
rect 2282 2679 2284 2687
rect 2287 2679 2289 2687
rect 2310 2685 2312 2693
rect 3120 2685 3122 2693
rect 2946 2672 2948 2680
rect 2962 2672 2964 2680
rect 2978 2672 2980 2680
rect 3001 2672 3003 2680
rect 3006 2672 3008 2680
rect 3032 2672 3034 2680
rect 3053 2672 3055 2680
rect 3073 2672 3075 2680
rect 3078 2672 3080 2680
rect 3096 2672 3098 2680
rect 3146 2679 3148 2687
rect 3151 2679 3153 2687
rect 3174 2685 3176 2693
rect 3201 2685 3203 2693
rect 3227 2679 3229 2687
rect 3232 2679 3234 2687
rect 3255 2685 3257 2693
rect 1635 2621 1637 2629
rect 1651 2621 1653 2629
rect 1656 2621 1658 2629
rect 1672 2621 1674 2629
rect 1688 2621 1690 2629
rect 1709 2621 1711 2629
rect 1714 2621 1716 2629
rect 1730 2621 1732 2629
rect 1746 2621 1748 2629
rect 1751 2621 1753 2629
rect 2580 2621 2582 2629
rect 2596 2621 2598 2629
rect 2601 2621 2603 2629
rect 2617 2621 2619 2629
rect 2633 2621 2635 2629
rect 2654 2621 2656 2629
rect 2659 2621 2661 2629
rect 2675 2621 2677 2629
rect 2691 2621 2693 2629
rect 2696 2621 2698 2629
rect 2001 2586 2003 2594
rect 2017 2586 2019 2594
rect 2033 2586 2035 2594
rect 2056 2586 2058 2594
rect 2061 2586 2063 2594
rect 2087 2586 2089 2594
rect 2108 2586 2110 2594
rect 2128 2586 2130 2594
rect 2133 2586 2135 2594
rect 2151 2586 2153 2594
rect 2201 2587 2203 2595
rect 2206 2587 2208 2595
rect 2282 2587 2284 2595
rect 2287 2587 2289 2595
rect 2946 2586 2948 2594
rect 2962 2586 2964 2594
rect 2978 2586 2980 2594
rect 3001 2586 3003 2594
rect 3006 2586 3008 2594
rect 3032 2586 3034 2594
rect 3053 2586 3055 2594
rect 3073 2586 3075 2594
rect 3078 2586 3080 2594
rect 3096 2586 3098 2594
rect 3146 2587 3148 2595
rect 3151 2587 3153 2595
rect 3227 2587 3229 2595
rect 3232 2587 3234 2595
rect 2001 2540 2003 2548
rect 2017 2540 2019 2548
rect 2033 2540 2035 2548
rect 2056 2540 2058 2548
rect 2061 2540 2063 2548
rect 2087 2540 2089 2548
rect 2108 2540 2110 2548
rect 2128 2540 2130 2548
rect 2133 2540 2135 2548
rect 2151 2540 2153 2548
rect 2201 2547 2203 2555
rect 2206 2547 2208 2555
rect 2229 2553 2231 2561
rect 2280 2553 2282 2561
rect 2306 2547 2308 2555
rect 2311 2547 2313 2555
rect 2334 2553 2336 2561
rect 2946 2540 2948 2548
rect 2962 2540 2964 2548
rect 2978 2540 2980 2548
rect 3001 2540 3003 2548
rect 3006 2540 3008 2548
rect 3032 2540 3034 2548
rect 3053 2540 3055 2548
rect 3073 2540 3075 2548
rect 3078 2540 3080 2548
rect 3096 2540 3098 2548
rect 3146 2547 3148 2555
rect 3151 2547 3153 2555
rect 3174 2553 3176 2561
rect 3225 2553 3227 2561
rect 3251 2547 3253 2555
rect 3256 2547 3258 2555
rect 3279 2553 3281 2561
rect 2001 2454 2003 2462
rect 2017 2454 2019 2462
rect 2033 2454 2035 2462
rect 2056 2454 2058 2462
rect 2061 2454 2063 2462
rect 2087 2454 2089 2462
rect 2108 2454 2110 2462
rect 2128 2454 2130 2462
rect 2133 2454 2135 2462
rect 2151 2454 2153 2462
rect 2201 2456 2203 2464
rect 2206 2456 2208 2464
rect 2306 2456 2308 2464
rect 2311 2456 2313 2464
rect 2946 2454 2948 2462
rect 2962 2454 2964 2462
rect 2978 2454 2980 2462
rect 3001 2454 3003 2462
rect 3006 2454 3008 2462
rect 3032 2454 3034 2462
rect 3053 2454 3055 2462
rect 3073 2454 3075 2462
rect 3078 2454 3080 2462
rect 3096 2454 3098 2462
rect 3146 2456 3148 2464
rect 3151 2456 3153 2464
rect 3251 2456 3253 2464
rect 3256 2456 3258 2464
rect 2001 2408 2003 2416
rect 2017 2408 2019 2416
rect 2033 2408 2035 2416
rect 2056 2408 2058 2416
rect 2061 2408 2063 2416
rect 2087 2408 2089 2416
rect 2108 2408 2110 2416
rect 2128 2408 2130 2416
rect 2133 2408 2135 2416
rect 2151 2408 2153 2416
rect 2201 2415 2203 2423
rect 2206 2415 2208 2423
rect 2229 2421 2231 2429
rect 2256 2421 2258 2429
rect 2282 2415 2284 2423
rect 2287 2415 2289 2423
rect 2310 2421 2312 2429
rect 2346 2421 2348 2429
rect 2372 2415 2374 2423
rect 2377 2415 2379 2423
rect 2400 2421 2402 2429
rect 2946 2408 2948 2416
rect 2962 2408 2964 2416
rect 2978 2408 2980 2416
rect 3001 2408 3003 2416
rect 3006 2408 3008 2416
rect 3032 2408 3034 2416
rect 3053 2408 3055 2416
rect 3073 2408 3075 2416
rect 3078 2408 3080 2416
rect 3096 2408 3098 2416
rect 3146 2415 3148 2423
rect 3151 2415 3153 2423
rect 3174 2421 3176 2429
rect 3201 2421 3203 2429
rect 3227 2415 3229 2423
rect 3232 2415 3234 2423
rect 3255 2421 3257 2429
rect 3291 2421 3293 2429
rect 3317 2415 3319 2423
rect 3322 2415 3324 2423
rect 3345 2421 3347 2429
rect 2001 2322 2003 2330
rect 2017 2322 2019 2330
rect 2033 2322 2035 2330
rect 2056 2322 2058 2330
rect 2061 2322 2063 2330
rect 2087 2322 2089 2330
rect 2108 2322 2110 2330
rect 2128 2322 2130 2330
rect 2133 2322 2135 2330
rect 2151 2322 2153 2330
rect 2201 2321 2203 2329
rect 2206 2321 2208 2329
rect 2282 2321 2284 2329
rect 2287 2321 2289 2329
rect 2372 2321 2374 2329
rect 2377 2321 2379 2329
rect 2946 2322 2948 2330
rect 2962 2322 2964 2330
rect 2978 2322 2980 2330
rect 3001 2322 3003 2330
rect 3006 2322 3008 2330
rect 3032 2322 3034 2330
rect 3053 2322 3055 2330
rect 3073 2322 3075 2330
rect 3078 2322 3080 2330
rect 3096 2322 3098 2330
rect 3146 2321 3148 2329
rect 3151 2321 3153 2329
rect 3227 2321 3229 2329
rect 3232 2321 3234 2329
rect 3317 2321 3319 2329
rect 3322 2321 3324 2329
rect 2001 2276 2003 2284
rect 2017 2276 2019 2284
rect 2033 2276 2035 2284
rect 2056 2276 2058 2284
rect 2061 2276 2063 2284
rect 2087 2276 2089 2284
rect 2108 2276 2110 2284
rect 2128 2276 2130 2284
rect 2133 2276 2135 2284
rect 2151 2276 2153 2284
rect 2201 2283 2203 2291
rect 2206 2283 2208 2291
rect 2229 2289 2231 2297
rect 2946 2276 2948 2284
rect 2962 2276 2964 2284
rect 2978 2276 2980 2284
rect 3001 2276 3003 2284
rect 3006 2276 3008 2284
rect 3032 2276 3034 2284
rect 3053 2276 3055 2284
rect 3073 2276 3075 2284
rect 3078 2276 3080 2284
rect 3096 2276 3098 2284
rect 3146 2283 3148 2291
rect 3151 2283 3153 2291
rect 3174 2289 3176 2297
rect 1512 2221 1514 2229
rect 1517 2221 1519 2229
rect 1533 2221 1535 2229
rect 1549 2221 1551 2229
rect 1554 2221 1556 2229
rect 1575 2221 1577 2229
rect 1591 2221 1593 2229
rect 1607 2221 1609 2229
rect 1612 2221 1614 2229
rect 1628 2221 1630 2229
rect 1644 2221 1646 2229
rect 1649 2221 1651 2229
rect 1665 2221 1667 2229
rect 1681 2221 1683 2229
rect 1686 2221 1688 2229
rect 1707 2221 1709 2229
rect 1723 2221 1725 2229
rect 1739 2221 1741 2229
rect 1744 2221 1746 2229
rect 1760 2221 1762 2229
rect 1776 2221 1778 2229
rect 1781 2221 1783 2229
rect 1797 2221 1799 2229
rect 1813 2221 1815 2229
rect 1818 2221 1820 2229
rect 1839 2221 1841 2229
rect 1855 2221 1857 2229
rect 1871 2221 1873 2229
rect 1876 2221 1878 2229
rect 1892 2221 1894 2229
rect 2457 2221 2459 2229
rect 2462 2221 2464 2229
rect 2478 2221 2480 2229
rect 2494 2221 2496 2229
rect 2499 2221 2501 2229
rect 2520 2221 2522 2229
rect 2536 2221 2538 2229
rect 2552 2221 2554 2229
rect 2557 2221 2559 2229
rect 2573 2221 2575 2229
rect 2589 2221 2591 2229
rect 2594 2221 2596 2229
rect 2610 2221 2612 2229
rect 2626 2221 2628 2229
rect 2631 2221 2633 2229
rect 2652 2221 2654 2229
rect 2668 2221 2670 2229
rect 2684 2221 2686 2229
rect 2689 2221 2691 2229
rect 2705 2221 2707 2229
rect 2721 2221 2723 2229
rect 2726 2221 2728 2229
rect 2742 2221 2744 2229
rect 2758 2221 2760 2229
rect 2763 2221 2765 2229
rect 2784 2221 2786 2229
rect 2800 2221 2802 2229
rect 2816 2221 2818 2229
rect 2821 2221 2823 2229
rect 2837 2221 2839 2229
rect 2001 2190 2003 2198
rect 2017 2190 2019 2198
rect 2033 2190 2035 2198
rect 2056 2190 2058 2198
rect 2061 2190 2063 2198
rect 2087 2190 2089 2198
rect 2108 2190 2110 2198
rect 2128 2190 2130 2198
rect 2133 2190 2135 2198
rect 2151 2190 2153 2198
rect 2201 2185 2203 2193
rect 2206 2185 2208 2193
rect 2235 2190 2237 2198
rect 2253 2190 2255 2198
rect 2278 2190 2280 2198
rect 2294 2190 2296 2198
rect 2317 2190 2319 2198
rect 2322 2190 2324 2198
rect 2348 2190 2350 2198
rect 2369 2190 2371 2198
rect 2389 2190 2391 2198
rect 2394 2190 2396 2198
rect 2412 2190 2414 2198
rect 2946 2190 2948 2198
rect 2962 2190 2964 2198
rect 2978 2190 2980 2198
rect 3001 2190 3003 2198
rect 3006 2190 3008 2198
rect 3032 2190 3034 2198
rect 3053 2190 3055 2198
rect 3073 2190 3075 2198
rect 3078 2190 3080 2198
rect 3096 2190 3098 2198
rect 3146 2185 3148 2193
rect 3151 2185 3153 2193
rect 3180 2190 3182 2198
rect 3198 2190 3200 2198
rect 3223 2190 3225 2198
rect 3239 2190 3241 2198
rect 3262 2190 3264 2198
rect 3267 2190 3269 2198
rect 3293 2190 3295 2198
rect 3314 2190 3316 2198
rect 3334 2190 3336 2198
rect 3339 2190 3341 2198
rect 3357 2190 3359 2198
rect 2295 2109 2297 2117
rect 2300 2109 2302 2117
rect 2316 2109 2318 2117
rect 2332 2109 2334 2117
rect 2337 2109 2339 2117
rect 2358 2109 2360 2117
rect 2374 2109 2376 2117
rect 2390 2109 2392 2117
rect 2395 2109 2397 2117
rect 2411 2109 2413 2117
rect 3240 2109 3242 2117
rect 3245 2109 3247 2117
rect 3261 2109 3263 2117
rect 3277 2109 3279 2117
rect 3282 2109 3284 2117
rect 3303 2109 3305 2117
rect 3319 2109 3321 2117
rect 3335 2109 3337 2117
rect 3340 2109 3342 2117
rect 3356 2109 3358 2117
rect 1512 2079 1514 2087
rect 1517 2079 1519 2087
rect 1533 2079 1535 2087
rect 1549 2079 1551 2087
rect 1554 2079 1556 2087
rect 1575 2079 1577 2087
rect 1591 2079 1593 2087
rect 1607 2079 1609 2087
rect 1612 2079 1614 2087
rect 1628 2079 1630 2087
rect 1644 2079 1646 2087
rect 1649 2079 1651 2087
rect 1665 2079 1667 2087
rect 1681 2079 1683 2087
rect 1686 2079 1688 2087
rect 1707 2079 1709 2087
rect 1723 2079 1725 2087
rect 1739 2079 1741 2087
rect 1744 2079 1746 2087
rect 1760 2079 1762 2087
rect 1776 2079 1778 2087
rect 1781 2079 1783 2087
rect 1797 2079 1799 2087
rect 1813 2079 1815 2087
rect 1818 2079 1820 2087
rect 1839 2079 1841 2087
rect 1855 2079 1857 2087
rect 1871 2079 1873 2087
rect 1876 2079 1878 2087
rect 1892 2079 1894 2087
rect 2457 2079 2459 2087
rect 2462 2079 2464 2087
rect 2478 2079 2480 2087
rect 2494 2079 2496 2087
rect 2499 2079 2501 2087
rect 2520 2079 2522 2087
rect 2536 2079 2538 2087
rect 2552 2079 2554 2087
rect 2557 2079 2559 2087
rect 2573 2079 2575 2087
rect 2589 2079 2591 2087
rect 2594 2079 2596 2087
rect 2610 2079 2612 2087
rect 2626 2079 2628 2087
rect 2631 2079 2633 2087
rect 2652 2079 2654 2087
rect 2668 2079 2670 2087
rect 2684 2079 2686 2087
rect 2689 2079 2691 2087
rect 2705 2079 2707 2087
rect 2721 2079 2723 2087
rect 2726 2079 2728 2087
rect 2742 2079 2744 2087
rect 2758 2079 2760 2087
rect 2763 2079 2765 2087
rect 2784 2079 2786 2087
rect 2800 2079 2802 2087
rect 2816 2079 2818 2087
rect 2821 2079 2823 2087
rect 2837 2079 2839 2087
rect 2295 2023 2297 2031
rect 2300 2023 2302 2031
rect 2316 2023 2318 2031
rect 2332 2023 2334 2031
rect 2337 2023 2339 2031
rect 2358 2023 2360 2031
rect 2374 2023 2376 2031
rect 2390 2023 2392 2031
rect 2395 2023 2397 2031
rect 2411 2023 2413 2031
rect 3240 2023 3242 2031
rect 3245 2023 3247 2031
rect 3261 2023 3263 2031
rect 3277 2023 3279 2031
rect 3282 2023 3284 2031
rect 3303 2023 3305 2031
rect 3319 2023 3321 2031
rect 3335 2023 3337 2031
rect 3340 2023 3342 2031
rect 3356 2023 3358 2031
rect 1512 1993 1514 2001
rect 1517 1993 1519 2001
rect 1533 1993 1535 2001
rect 1549 1993 1551 2001
rect 1554 1993 1556 2001
rect 1575 1993 1577 2001
rect 1591 1993 1593 2001
rect 1607 1993 1609 2001
rect 1612 1993 1614 2001
rect 1628 1993 1630 2001
rect 1644 1993 1646 2001
rect 1649 1993 1651 2001
rect 1665 1993 1667 2001
rect 1681 1993 1683 2001
rect 1686 1993 1688 2001
rect 1707 1993 1709 2001
rect 1723 1993 1725 2001
rect 1739 1993 1741 2001
rect 1744 1993 1746 2001
rect 1760 1993 1762 2001
rect 1776 1993 1778 2001
rect 1781 1993 1783 2001
rect 1797 1993 1799 2001
rect 1813 1993 1815 2001
rect 1818 1993 1820 2001
rect 1839 1993 1841 2001
rect 1855 1993 1857 2001
rect 1871 1993 1873 2001
rect 1876 1993 1878 2001
rect 1892 1993 1894 2001
rect 2457 1993 2459 2001
rect 2462 1993 2464 2001
rect 2478 1993 2480 2001
rect 2494 1993 2496 2001
rect 2499 1993 2501 2001
rect 2520 1993 2522 2001
rect 2536 1993 2538 2001
rect 2552 1993 2554 2001
rect 2557 1993 2559 2001
rect 2573 1993 2575 2001
rect 2589 1993 2591 2001
rect 2594 1993 2596 2001
rect 2610 1993 2612 2001
rect 2626 1993 2628 2001
rect 2631 1993 2633 2001
rect 2652 1993 2654 2001
rect 2668 1993 2670 2001
rect 2684 1993 2686 2001
rect 2689 1993 2691 2001
rect 2705 1993 2707 2001
rect 2721 1993 2723 2001
rect 2726 1993 2728 2001
rect 2742 1993 2744 2001
rect 2758 1993 2760 2001
rect 2763 1993 2765 2001
rect 2784 1993 2786 2001
rect 2800 1993 2802 2001
rect 2816 1993 2818 2001
rect 2821 1993 2823 2001
rect 2837 1993 2839 2001
rect 1512 1853 1514 1861
rect 1517 1853 1519 1861
rect 1533 1853 1535 1861
rect 1549 1853 1551 1861
rect 1554 1853 1556 1861
rect 1575 1853 1577 1861
rect 1591 1853 1593 1861
rect 1607 1853 1609 1861
rect 1612 1853 1614 1861
rect 1628 1853 1630 1861
rect 1644 1853 1646 1861
rect 1649 1853 1651 1861
rect 1665 1853 1667 1861
rect 1681 1853 1683 1861
rect 1686 1853 1688 1861
rect 1707 1853 1709 1861
rect 1723 1853 1725 1861
rect 1739 1853 1741 1861
rect 1744 1853 1746 1861
rect 1760 1853 1762 1861
rect 1776 1853 1778 1861
rect 1781 1853 1783 1861
rect 1797 1853 1799 1861
rect 1813 1853 1815 1861
rect 1818 1853 1820 1861
rect 1839 1853 1841 1861
rect 1855 1853 1857 1861
rect 1871 1853 1873 1861
rect 1876 1853 1878 1861
rect 1892 1853 1894 1861
rect 2457 1853 2459 1861
rect 2462 1853 2464 1861
rect 2478 1853 2480 1861
rect 2494 1853 2496 1861
rect 2499 1853 2501 1861
rect 2520 1853 2522 1861
rect 2536 1853 2538 1861
rect 2552 1853 2554 1861
rect 2557 1853 2559 1861
rect 2573 1853 2575 1861
rect 2589 1853 2591 1861
rect 2594 1853 2596 1861
rect 2610 1853 2612 1861
rect 2626 1853 2628 1861
rect 2631 1853 2633 1861
rect 2652 1853 2654 1861
rect 2668 1853 2670 1861
rect 2684 1853 2686 1861
rect 2689 1853 2691 1861
rect 2705 1853 2707 1861
rect 2721 1853 2723 1861
rect 2726 1853 2728 1861
rect 2742 1853 2744 1861
rect 2758 1853 2760 1861
rect 2763 1853 2765 1861
rect 2784 1853 2786 1861
rect 2800 1853 2802 1861
rect 2816 1853 2818 1861
rect 2821 1853 2823 1861
rect 2837 1853 2839 1861
<< ndiffusion >>
rect 2700 4250 2701 4254
rect 2703 4250 2704 4254
rect 2724 4246 2727 4250
rect 2729 4246 2732 4250
rect 2734 4246 2735 4250
rect 2754 4242 2755 4246
rect 2757 4242 2758 4246
rect 2886 4211 2887 4223
rect 2889 4211 2890 4223
rect 2939 4211 2940 4223
rect 2942 4211 2943 4223
rect 2724 4186 2727 4190
rect 2729 4186 2732 4190
rect 2734 4186 2735 4190
rect 2678 4120 2679 4124
rect 2681 4120 2682 4124
rect 2700 4120 2701 4124
rect 2703 4120 2704 4124
rect 2724 4116 2727 4120
rect 2729 4116 2732 4120
rect 2734 4116 2735 4120
rect 2754 4112 2755 4116
rect 2757 4112 2758 4116
rect 2792 4081 2793 4093
rect 2795 4081 2796 4093
rect 2845 4081 2846 4093
rect 2848 4081 2849 4093
rect 2724 4056 2727 4060
rect 2729 4056 2732 4060
rect 2734 4056 2735 4060
rect 1995 3715 1996 3719
rect 1998 3715 2001 3719
rect 2003 3715 2004 3719
rect 2016 3715 2017 3719
rect 2019 3715 2020 3719
rect 2032 3715 2033 3719
rect 2035 3715 2038 3719
rect 2040 3715 2041 3719
rect 2058 3715 2059 3719
rect 2061 3715 2062 3719
rect 2074 3715 2075 3719
rect 2077 3715 2078 3719
rect 2090 3715 2091 3719
rect 2093 3715 2096 3719
rect 2098 3715 2099 3719
rect 2111 3715 2112 3719
rect 2114 3715 2115 3719
rect 2127 3715 2128 3719
rect 2130 3715 2133 3719
rect 2135 3715 2136 3719
rect 2148 3715 2149 3719
rect 2151 3715 2152 3719
rect 2164 3715 2165 3719
rect 2167 3715 2170 3719
rect 2172 3715 2173 3719
rect 2190 3715 2191 3719
rect 2193 3715 2194 3719
rect 2206 3715 2207 3719
rect 2209 3715 2210 3719
rect 2222 3715 2223 3719
rect 2225 3715 2228 3719
rect 2230 3715 2231 3719
rect 2243 3715 2244 3719
rect 2246 3715 2247 3719
rect 2259 3715 2260 3719
rect 2262 3715 2265 3719
rect 2267 3715 2268 3719
rect 2280 3715 2281 3719
rect 2283 3715 2284 3719
rect 2296 3715 2297 3719
rect 2299 3715 2302 3719
rect 2304 3715 2305 3719
rect 2322 3715 2323 3719
rect 2325 3715 2326 3719
rect 2338 3715 2339 3719
rect 2341 3715 2342 3719
rect 2354 3715 2355 3719
rect 2357 3715 2360 3719
rect 2362 3715 2363 3719
rect 2375 3715 2376 3719
rect 2378 3715 2379 3719
rect 2391 3715 2392 3719
rect 2394 3715 2397 3719
rect 2399 3715 2400 3719
rect 2412 3715 2413 3719
rect 2415 3715 2416 3719
rect 2428 3715 2429 3719
rect 2431 3715 2434 3719
rect 2436 3715 2437 3719
rect 2454 3715 2455 3719
rect 2457 3715 2458 3719
rect 2470 3715 2471 3719
rect 2473 3715 2474 3719
rect 2486 3715 2487 3719
rect 2489 3715 2492 3719
rect 2494 3715 2495 3719
rect 2507 3715 2508 3719
rect 2510 3715 2511 3719
rect 2940 3715 2941 3719
rect 2943 3715 2946 3719
rect 2948 3715 2949 3719
rect 2961 3715 2962 3719
rect 2964 3715 2965 3719
rect 2977 3715 2978 3719
rect 2980 3715 2983 3719
rect 2985 3715 2986 3719
rect 3003 3715 3004 3719
rect 3006 3715 3007 3719
rect 3019 3715 3020 3719
rect 3022 3715 3023 3719
rect 3035 3715 3036 3719
rect 3038 3715 3041 3719
rect 3043 3715 3044 3719
rect 3056 3715 3057 3719
rect 3059 3715 3060 3719
rect 3072 3715 3073 3719
rect 3075 3715 3078 3719
rect 3080 3715 3081 3719
rect 3093 3715 3094 3719
rect 3096 3715 3097 3719
rect 3109 3715 3110 3719
rect 3112 3715 3115 3719
rect 3117 3715 3118 3719
rect 3135 3715 3136 3719
rect 3138 3715 3139 3719
rect 3151 3715 3152 3719
rect 3154 3715 3155 3719
rect 3167 3715 3168 3719
rect 3170 3715 3173 3719
rect 3175 3715 3176 3719
rect 3188 3715 3189 3719
rect 3191 3715 3192 3719
rect 3204 3715 3205 3719
rect 3207 3715 3210 3719
rect 3212 3715 3213 3719
rect 3225 3715 3226 3719
rect 3228 3715 3229 3719
rect 3241 3715 3242 3719
rect 3244 3715 3247 3719
rect 3249 3715 3250 3719
rect 3267 3715 3268 3719
rect 3270 3715 3271 3719
rect 3283 3715 3284 3719
rect 3286 3715 3287 3719
rect 3299 3715 3300 3719
rect 3302 3715 3305 3719
rect 3307 3715 3308 3719
rect 3320 3715 3321 3719
rect 3323 3715 3324 3719
rect 3336 3715 3337 3719
rect 3339 3715 3342 3719
rect 3344 3715 3345 3719
rect 3357 3715 3358 3719
rect 3360 3715 3361 3719
rect 3373 3715 3374 3719
rect 3376 3715 3379 3719
rect 3381 3715 3382 3719
rect 3399 3715 3400 3719
rect 3402 3715 3403 3719
rect 3415 3715 3416 3719
rect 3418 3715 3419 3719
rect 3431 3715 3432 3719
rect 3434 3715 3437 3719
rect 3439 3715 3440 3719
rect 3452 3715 3453 3719
rect 3455 3715 3456 3719
rect 1643 3682 1644 3686
rect 1646 3682 1649 3686
rect 1651 3682 1652 3686
rect 1664 3682 1665 3686
rect 1667 3682 1668 3686
rect 1680 3682 1681 3686
rect 1683 3682 1686 3686
rect 1688 3682 1689 3686
rect 1706 3682 1707 3686
rect 1709 3682 1710 3686
rect 1722 3682 1723 3686
rect 1725 3682 1726 3686
rect 1738 3682 1739 3686
rect 1741 3682 1744 3686
rect 1746 3682 1747 3686
rect 1759 3682 1760 3686
rect 1762 3682 1763 3686
rect 2588 3682 2589 3686
rect 2591 3682 2594 3686
rect 2596 3682 2597 3686
rect 2609 3682 2610 3686
rect 2612 3682 2613 3686
rect 2625 3682 2626 3686
rect 2628 3682 2631 3686
rect 2633 3682 2634 3686
rect 2651 3682 2652 3686
rect 2654 3682 2655 3686
rect 2667 3682 2668 3686
rect 2670 3682 2671 3686
rect 2683 3682 2684 3686
rect 2686 3682 2689 3686
rect 2691 3682 2692 3686
rect 2704 3682 2705 3686
rect 2707 3682 2708 3686
rect 1767 3645 1768 3649
rect 1770 3645 1771 3649
rect 2174 3649 2175 3653
rect 2177 3649 2178 3653
rect 2198 3645 2201 3649
rect 2203 3645 2206 3649
rect 2208 3645 2209 3649
rect 2255 3649 2256 3653
rect 2258 3649 2259 3653
rect 2279 3645 2282 3649
rect 2284 3645 2287 3649
rect 2289 3645 2290 3649
rect 2228 3641 2229 3645
rect 2231 3641 2232 3645
rect 1650 3636 1651 3640
rect 1653 3636 1654 3640
rect 2000 3636 2001 3640
rect 2003 3636 2004 3640
rect 2016 3636 2017 3640
rect 2019 3636 2020 3640
rect 2032 3636 2033 3640
rect 2035 3636 2036 3640
rect 2051 3636 2056 3640
rect 2058 3636 2061 3640
rect 2063 3636 2064 3640
rect 2085 3636 2087 3640
rect 2089 3636 2090 3640
rect 2107 3636 2108 3640
rect 2110 3636 2111 3640
rect 2123 3636 2128 3640
rect 2130 3636 2133 3640
rect 2135 3636 2136 3640
rect 2150 3636 2151 3640
rect 2153 3636 2154 3640
rect 2309 3641 2310 3645
rect 2312 3641 2313 3645
rect 2712 3645 2713 3649
rect 2715 3645 2716 3649
rect 3119 3649 3120 3653
rect 3122 3649 3123 3653
rect 3143 3645 3146 3649
rect 3148 3645 3151 3649
rect 3153 3645 3154 3649
rect 3200 3649 3201 3653
rect 3203 3649 3204 3653
rect 3224 3645 3227 3649
rect 3229 3645 3232 3649
rect 3234 3645 3235 3649
rect 3173 3641 3174 3645
rect 3176 3641 3177 3645
rect 2595 3636 2596 3640
rect 2598 3636 2599 3640
rect 2945 3636 2946 3640
rect 2948 3636 2949 3640
rect 2961 3636 2962 3640
rect 2964 3636 2965 3640
rect 2977 3636 2978 3640
rect 2980 3636 2981 3640
rect 2996 3636 3001 3640
rect 3003 3636 3006 3640
rect 3008 3636 3009 3640
rect 3030 3636 3032 3640
rect 3034 3636 3035 3640
rect 3052 3636 3053 3640
rect 3055 3636 3056 3640
rect 3068 3636 3073 3640
rect 3075 3636 3078 3640
rect 3080 3636 3081 3640
rect 3095 3636 3096 3640
rect 3098 3636 3099 3640
rect 3254 3641 3255 3645
rect 3257 3641 3258 3645
rect 2000 3590 2001 3594
rect 2003 3590 2004 3594
rect 2016 3590 2017 3594
rect 2019 3590 2020 3594
rect 2032 3590 2033 3594
rect 2035 3590 2036 3594
rect 2051 3590 2056 3594
rect 2058 3590 2061 3594
rect 2063 3590 2064 3594
rect 2085 3590 2087 3594
rect 2089 3590 2090 3594
rect 2107 3590 2108 3594
rect 2110 3590 2111 3594
rect 2123 3590 2128 3594
rect 2130 3590 2133 3594
rect 2135 3590 2136 3594
rect 2150 3590 2151 3594
rect 2153 3590 2154 3594
rect 1634 3580 1635 3584
rect 1637 3580 1638 3584
rect 1650 3580 1651 3584
rect 1653 3580 1656 3584
rect 1658 3580 1659 3584
rect 1671 3580 1672 3584
rect 1674 3580 1675 3584
rect 1687 3580 1688 3584
rect 1690 3580 1691 3584
rect 1708 3580 1709 3584
rect 1711 3580 1714 3584
rect 1716 3580 1717 3584
rect 1729 3580 1730 3584
rect 1732 3580 1733 3584
rect 1745 3580 1746 3584
rect 1748 3580 1751 3584
rect 1753 3580 1754 3584
rect 2198 3589 2201 3593
rect 2203 3589 2206 3593
rect 2208 3589 2209 3593
rect 2279 3589 2282 3593
rect 2284 3589 2287 3593
rect 2289 3589 2290 3593
rect 2945 3590 2946 3594
rect 2948 3590 2949 3594
rect 2961 3590 2962 3594
rect 2964 3590 2965 3594
rect 2977 3590 2978 3594
rect 2980 3590 2981 3594
rect 2996 3590 3001 3594
rect 3003 3590 3006 3594
rect 3008 3590 3009 3594
rect 3030 3590 3032 3594
rect 3034 3590 3035 3594
rect 3052 3590 3053 3594
rect 3055 3590 3056 3594
rect 3068 3590 3073 3594
rect 3075 3590 3078 3594
rect 3080 3590 3081 3594
rect 3095 3590 3096 3594
rect 3098 3590 3099 3594
rect 2579 3580 2580 3584
rect 2582 3580 2583 3584
rect 2595 3580 2596 3584
rect 2598 3580 2601 3584
rect 2603 3580 2604 3584
rect 2616 3580 2617 3584
rect 2619 3580 2620 3584
rect 2632 3580 2633 3584
rect 2635 3580 2636 3584
rect 2653 3580 2654 3584
rect 2656 3580 2659 3584
rect 2661 3580 2662 3584
rect 2674 3580 2675 3584
rect 2677 3580 2678 3584
rect 2690 3580 2691 3584
rect 2693 3580 2696 3584
rect 2698 3580 2699 3584
rect 3143 3589 3146 3593
rect 3148 3589 3151 3593
rect 3153 3589 3154 3593
rect 3224 3589 3227 3593
rect 3229 3589 3232 3593
rect 3234 3589 3235 3593
rect 2198 3513 2201 3517
rect 2203 3513 2206 3517
rect 2208 3513 2209 3517
rect 2279 3517 2280 3521
rect 2282 3517 2283 3521
rect 2303 3513 2306 3517
rect 2308 3513 2311 3517
rect 2313 3513 2314 3517
rect 2228 3509 2229 3513
rect 2231 3509 2232 3513
rect 2000 3504 2001 3508
rect 2003 3504 2004 3508
rect 2016 3504 2017 3508
rect 2019 3504 2020 3508
rect 2032 3504 2033 3508
rect 2035 3504 2036 3508
rect 2051 3504 2056 3508
rect 2058 3504 2061 3508
rect 2063 3504 2064 3508
rect 2085 3504 2087 3508
rect 2089 3504 2090 3508
rect 2107 3504 2108 3508
rect 2110 3504 2111 3508
rect 2123 3504 2128 3508
rect 2130 3504 2133 3508
rect 2135 3504 2136 3508
rect 2150 3504 2151 3508
rect 2153 3504 2154 3508
rect 2333 3509 2334 3513
rect 2336 3509 2337 3513
rect 3143 3513 3146 3517
rect 3148 3513 3151 3517
rect 3153 3513 3154 3517
rect 3224 3517 3225 3521
rect 3227 3517 3228 3521
rect 3248 3513 3251 3517
rect 3253 3513 3256 3517
rect 3258 3513 3259 3517
rect 3173 3509 3174 3513
rect 3176 3509 3177 3513
rect 2945 3504 2946 3508
rect 2948 3504 2949 3508
rect 2961 3504 2962 3508
rect 2964 3504 2965 3508
rect 2977 3504 2978 3508
rect 2980 3504 2981 3508
rect 2996 3504 3001 3508
rect 3003 3504 3006 3508
rect 3008 3504 3009 3508
rect 3030 3504 3032 3508
rect 3034 3504 3035 3508
rect 3052 3504 3053 3508
rect 3055 3504 3056 3508
rect 3068 3504 3073 3508
rect 3075 3504 3078 3508
rect 3080 3504 3081 3508
rect 3095 3504 3096 3508
rect 3098 3504 3099 3508
rect 3278 3509 3279 3513
rect 3281 3509 3282 3513
rect 2000 3458 2001 3462
rect 2003 3458 2004 3462
rect 2016 3458 2017 3462
rect 2019 3458 2020 3462
rect 2032 3458 2033 3462
rect 2035 3458 2036 3462
rect 2051 3458 2056 3462
rect 2058 3458 2061 3462
rect 2063 3458 2064 3462
rect 2085 3458 2087 3462
rect 2089 3458 2090 3462
rect 2107 3458 2108 3462
rect 2110 3458 2111 3462
rect 2123 3458 2128 3462
rect 2130 3458 2133 3462
rect 2135 3458 2136 3462
rect 2150 3458 2151 3462
rect 2153 3458 2154 3462
rect 2198 3458 2201 3462
rect 2203 3458 2206 3462
rect 2208 3458 2209 3462
rect 2303 3458 2306 3462
rect 2308 3458 2311 3462
rect 2313 3458 2314 3462
rect 2945 3458 2946 3462
rect 2948 3458 2949 3462
rect 2961 3458 2962 3462
rect 2964 3458 2965 3462
rect 2977 3458 2978 3462
rect 2980 3458 2981 3462
rect 2996 3458 3001 3462
rect 3003 3458 3006 3462
rect 3008 3458 3009 3462
rect 3030 3458 3032 3462
rect 3034 3458 3035 3462
rect 3052 3458 3053 3462
rect 3055 3458 3056 3462
rect 3068 3458 3073 3462
rect 3075 3458 3078 3462
rect 3080 3458 3081 3462
rect 3095 3458 3096 3462
rect 3098 3458 3099 3462
rect 3143 3458 3146 3462
rect 3148 3458 3151 3462
rect 3153 3458 3154 3462
rect 3248 3458 3251 3462
rect 3253 3458 3256 3462
rect 3258 3458 3259 3462
rect 2198 3381 2201 3385
rect 2203 3381 2206 3385
rect 2208 3381 2209 3385
rect 2255 3385 2256 3389
rect 2258 3385 2259 3389
rect 2279 3381 2282 3385
rect 2284 3381 2287 3385
rect 2289 3381 2290 3385
rect 2345 3385 2346 3389
rect 2348 3385 2349 3389
rect 2369 3381 2372 3385
rect 2374 3381 2377 3385
rect 2379 3381 2380 3385
rect 2228 3377 2229 3381
rect 2231 3377 2232 3381
rect 2000 3372 2001 3376
rect 2003 3372 2004 3376
rect 2016 3372 2017 3376
rect 2019 3372 2020 3376
rect 2032 3372 2033 3376
rect 2035 3372 2036 3376
rect 2051 3372 2056 3376
rect 2058 3372 2061 3376
rect 2063 3372 2064 3376
rect 2085 3372 2087 3376
rect 2089 3372 2090 3376
rect 2107 3372 2108 3376
rect 2110 3372 2111 3376
rect 2123 3372 2128 3376
rect 2130 3372 2133 3376
rect 2135 3372 2136 3376
rect 2150 3372 2151 3376
rect 2153 3372 2154 3376
rect 2309 3377 2310 3381
rect 2312 3377 2313 3381
rect 2399 3377 2400 3381
rect 2402 3377 2403 3381
rect 3143 3381 3146 3385
rect 3148 3381 3151 3385
rect 3153 3381 3154 3385
rect 3200 3385 3201 3389
rect 3203 3385 3204 3389
rect 3224 3381 3227 3385
rect 3229 3381 3232 3385
rect 3234 3381 3235 3385
rect 3290 3385 3291 3389
rect 3293 3385 3294 3389
rect 3314 3381 3317 3385
rect 3319 3381 3322 3385
rect 3324 3381 3325 3385
rect 3173 3377 3174 3381
rect 3176 3377 3177 3381
rect 2945 3372 2946 3376
rect 2948 3372 2949 3376
rect 2961 3372 2962 3376
rect 2964 3372 2965 3376
rect 2977 3372 2978 3376
rect 2980 3372 2981 3376
rect 2996 3372 3001 3376
rect 3003 3372 3006 3376
rect 3008 3372 3009 3376
rect 3030 3372 3032 3376
rect 3034 3372 3035 3376
rect 3052 3372 3053 3376
rect 3055 3372 3056 3376
rect 3068 3372 3073 3376
rect 3075 3372 3078 3376
rect 3080 3372 3081 3376
rect 3095 3372 3096 3376
rect 3098 3372 3099 3376
rect 3254 3377 3255 3381
rect 3257 3377 3258 3381
rect 3344 3377 3345 3381
rect 3347 3377 3348 3381
rect 2000 3326 2001 3330
rect 2003 3326 2004 3330
rect 2016 3326 2017 3330
rect 2019 3326 2020 3330
rect 2032 3326 2033 3330
rect 2035 3326 2036 3330
rect 2051 3326 2056 3330
rect 2058 3326 2061 3330
rect 2063 3326 2064 3330
rect 2085 3326 2087 3330
rect 2089 3326 2090 3330
rect 2107 3326 2108 3330
rect 2110 3326 2111 3330
rect 2123 3326 2128 3330
rect 2130 3326 2133 3330
rect 2135 3326 2136 3330
rect 2150 3326 2151 3330
rect 2153 3326 2154 3330
rect 2198 3323 2201 3327
rect 2203 3323 2206 3327
rect 2208 3323 2209 3327
rect 2279 3323 2282 3327
rect 2284 3323 2287 3327
rect 2289 3323 2290 3327
rect 2369 3323 2372 3327
rect 2374 3323 2377 3327
rect 2379 3323 2380 3327
rect 2945 3326 2946 3330
rect 2948 3326 2949 3330
rect 2961 3326 2962 3330
rect 2964 3326 2965 3330
rect 2977 3326 2978 3330
rect 2980 3326 2981 3330
rect 2996 3326 3001 3330
rect 3003 3326 3006 3330
rect 3008 3326 3009 3330
rect 3030 3326 3032 3330
rect 3034 3326 3035 3330
rect 3052 3326 3053 3330
rect 3055 3326 3056 3330
rect 3068 3326 3073 3330
rect 3075 3326 3078 3330
rect 3080 3326 3081 3330
rect 3095 3326 3096 3330
rect 3098 3326 3099 3330
rect 3143 3323 3146 3327
rect 3148 3323 3151 3327
rect 3153 3323 3154 3327
rect 3224 3323 3227 3327
rect 3229 3323 3232 3327
rect 3234 3323 3235 3327
rect 3314 3323 3317 3327
rect 3319 3323 3322 3327
rect 3324 3323 3325 3327
rect 2198 3249 2201 3253
rect 2203 3249 2206 3253
rect 2208 3249 2209 3253
rect 2228 3245 2229 3249
rect 2231 3245 2232 3249
rect 2000 3240 2001 3244
rect 2003 3240 2004 3244
rect 2016 3240 2017 3244
rect 2019 3240 2020 3244
rect 2032 3240 2033 3244
rect 2035 3240 2036 3244
rect 2051 3240 2056 3244
rect 2058 3240 2061 3244
rect 2063 3240 2064 3244
rect 2085 3240 2087 3244
rect 2089 3240 2090 3244
rect 2107 3240 2108 3244
rect 2110 3240 2111 3244
rect 2123 3240 2128 3244
rect 2130 3240 2133 3244
rect 2135 3240 2136 3244
rect 2150 3240 2151 3244
rect 2153 3240 2154 3244
rect 3143 3249 3146 3253
rect 3148 3249 3151 3253
rect 3153 3249 3154 3253
rect 3173 3245 3174 3249
rect 3176 3245 3177 3249
rect 2945 3240 2946 3244
rect 2948 3240 2949 3244
rect 2961 3240 2962 3244
rect 2964 3240 2965 3244
rect 2977 3240 2978 3244
rect 2980 3240 2981 3244
rect 2996 3240 3001 3244
rect 3003 3240 3006 3244
rect 3008 3240 3009 3244
rect 3030 3240 3032 3244
rect 3034 3240 3035 3244
rect 3052 3240 3053 3244
rect 3055 3240 3056 3244
rect 3068 3240 3073 3244
rect 3075 3240 3078 3244
rect 3080 3240 3081 3244
rect 3095 3240 3096 3244
rect 3098 3240 3099 3244
rect 2000 3194 2001 3198
rect 2003 3194 2004 3198
rect 2016 3194 2017 3198
rect 2019 3194 2020 3198
rect 2032 3194 2033 3198
rect 2035 3194 2036 3198
rect 2051 3194 2056 3198
rect 2058 3194 2061 3198
rect 2063 3194 2064 3198
rect 2085 3194 2087 3198
rect 2089 3194 2090 3198
rect 2107 3194 2108 3198
rect 2110 3194 2111 3198
rect 2123 3194 2128 3198
rect 2130 3194 2133 3198
rect 2135 3194 2136 3198
rect 2150 3194 2151 3198
rect 2153 3194 2154 3198
rect 2234 3194 2235 3198
rect 2237 3194 2238 3198
rect 2242 3194 2248 3198
rect 2252 3194 2253 3198
rect 2255 3194 2256 3198
rect 2277 3194 2278 3198
rect 2280 3194 2281 3198
rect 2293 3194 2294 3198
rect 2296 3194 2297 3198
rect 2312 3194 2317 3198
rect 2319 3194 2322 3198
rect 2324 3194 2325 3198
rect 2346 3194 2348 3198
rect 2350 3194 2351 3198
rect 2368 3194 2369 3198
rect 2371 3194 2372 3198
rect 2384 3194 2389 3198
rect 2391 3194 2394 3198
rect 2396 3194 2397 3198
rect 2411 3194 2412 3198
rect 2414 3194 2415 3198
rect 1511 3180 1512 3184
rect 1514 3180 1517 3184
rect 1519 3180 1520 3184
rect 1532 3180 1533 3184
rect 1535 3180 1536 3184
rect 1548 3180 1549 3184
rect 1551 3180 1554 3184
rect 1556 3180 1557 3184
rect 1574 3180 1575 3184
rect 1577 3180 1578 3184
rect 1590 3180 1591 3184
rect 1593 3180 1594 3184
rect 1606 3180 1607 3184
rect 1609 3180 1612 3184
rect 1614 3180 1615 3184
rect 1627 3180 1628 3184
rect 1630 3180 1631 3184
rect 1643 3180 1644 3184
rect 1646 3180 1649 3184
rect 1651 3180 1652 3184
rect 1664 3180 1665 3184
rect 1667 3180 1668 3184
rect 1680 3180 1681 3184
rect 1683 3180 1686 3184
rect 1688 3180 1689 3184
rect 1706 3180 1707 3184
rect 1709 3180 1710 3184
rect 1722 3180 1723 3184
rect 1725 3180 1726 3184
rect 1738 3180 1739 3184
rect 1741 3180 1744 3184
rect 1746 3180 1747 3184
rect 1759 3180 1760 3184
rect 1762 3180 1763 3184
rect 1775 3180 1776 3184
rect 1778 3180 1781 3184
rect 1783 3180 1784 3184
rect 1796 3180 1797 3184
rect 1799 3180 1800 3184
rect 1812 3180 1813 3184
rect 1815 3180 1818 3184
rect 1820 3180 1821 3184
rect 1838 3180 1839 3184
rect 1841 3180 1842 3184
rect 1854 3180 1855 3184
rect 1857 3180 1858 3184
rect 1870 3180 1871 3184
rect 1873 3180 1876 3184
rect 1878 3180 1879 3184
rect 1891 3180 1892 3184
rect 1894 3180 1895 3184
rect 2198 3187 2201 3191
rect 2203 3187 2206 3191
rect 2208 3187 2209 3191
rect 2945 3194 2946 3198
rect 2948 3194 2949 3198
rect 2961 3194 2962 3198
rect 2964 3194 2965 3198
rect 2977 3194 2978 3198
rect 2980 3194 2981 3198
rect 2996 3194 3001 3198
rect 3003 3194 3006 3198
rect 3008 3194 3009 3198
rect 3030 3194 3032 3198
rect 3034 3194 3035 3198
rect 3052 3194 3053 3198
rect 3055 3194 3056 3198
rect 3068 3194 3073 3198
rect 3075 3194 3078 3198
rect 3080 3194 3081 3198
rect 3095 3194 3096 3198
rect 3098 3194 3099 3198
rect 3179 3194 3180 3198
rect 3182 3194 3183 3198
rect 3187 3194 3193 3198
rect 3197 3194 3198 3198
rect 3200 3194 3201 3198
rect 3222 3194 3223 3198
rect 3225 3194 3226 3198
rect 3238 3194 3239 3198
rect 3241 3194 3242 3198
rect 3257 3194 3262 3198
rect 3264 3194 3267 3198
rect 3269 3194 3270 3198
rect 3291 3194 3293 3198
rect 3295 3194 3296 3198
rect 3313 3194 3314 3198
rect 3316 3194 3317 3198
rect 3329 3194 3334 3198
rect 3336 3194 3339 3198
rect 3341 3194 3342 3198
rect 3356 3194 3357 3198
rect 3359 3194 3360 3198
rect 2456 3180 2457 3184
rect 2459 3180 2462 3184
rect 2464 3180 2465 3184
rect 2477 3180 2478 3184
rect 2480 3180 2481 3184
rect 2493 3180 2494 3184
rect 2496 3180 2499 3184
rect 2501 3180 2502 3184
rect 2519 3180 2520 3184
rect 2522 3180 2523 3184
rect 2535 3180 2536 3184
rect 2538 3180 2539 3184
rect 2551 3180 2552 3184
rect 2554 3180 2557 3184
rect 2559 3180 2560 3184
rect 2572 3180 2573 3184
rect 2575 3180 2576 3184
rect 2588 3180 2589 3184
rect 2591 3180 2594 3184
rect 2596 3180 2597 3184
rect 2609 3180 2610 3184
rect 2612 3180 2613 3184
rect 2625 3180 2626 3184
rect 2628 3180 2631 3184
rect 2633 3180 2634 3184
rect 2651 3180 2652 3184
rect 2654 3180 2655 3184
rect 2667 3180 2668 3184
rect 2670 3180 2671 3184
rect 2683 3180 2684 3184
rect 2686 3180 2689 3184
rect 2691 3180 2692 3184
rect 2704 3180 2705 3184
rect 2707 3180 2708 3184
rect 2720 3180 2721 3184
rect 2723 3180 2726 3184
rect 2728 3180 2729 3184
rect 2741 3180 2742 3184
rect 2744 3180 2745 3184
rect 2757 3180 2758 3184
rect 2760 3180 2763 3184
rect 2765 3180 2766 3184
rect 2783 3180 2784 3184
rect 2786 3180 2787 3184
rect 2799 3180 2800 3184
rect 2802 3180 2803 3184
rect 2815 3180 2816 3184
rect 2818 3180 2821 3184
rect 2823 3180 2824 3184
rect 2836 3180 2837 3184
rect 2839 3180 2840 3184
rect 3143 3187 3146 3191
rect 3148 3187 3151 3191
rect 3153 3187 3154 3191
rect 1626 3136 1627 3140
rect 1629 3136 1630 3140
rect 1650 3136 1651 3140
rect 1653 3136 1654 3140
rect 2424 3140 2428 3141
rect 2424 3137 2428 3138
rect 2571 3136 2572 3140
rect 2574 3136 2575 3140
rect 2595 3136 2596 3140
rect 2598 3136 2599 3140
rect 3369 3140 3373 3141
rect 3369 3137 3373 3138
rect 1646 3123 1647 3127
rect 1649 3123 1650 3127
rect 2591 3123 2592 3127
rect 2594 3123 2595 3127
rect 1638 3111 1642 3112
rect 1638 3108 1642 3109
rect 2583 3111 2587 3112
rect 2583 3108 2587 3109
rect 1626 3100 1627 3104
rect 1629 3100 1630 3104
rect 1650 3100 1651 3104
rect 1653 3100 1654 3104
rect 2571 3100 2572 3104
rect 2574 3100 2575 3104
rect 2595 3100 2596 3104
rect 2598 3100 2599 3104
rect 2294 3068 2295 3072
rect 2297 3068 2300 3072
rect 2302 3068 2303 3072
rect 2315 3068 2316 3072
rect 2318 3068 2319 3072
rect 2331 3068 2332 3072
rect 2334 3068 2337 3072
rect 2339 3068 2340 3072
rect 2357 3068 2358 3072
rect 2360 3068 2361 3072
rect 2373 3068 2374 3072
rect 2376 3068 2377 3072
rect 2389 3068 2390 3072
rect 2392 3068 2395 3072
rect 2397 3068 2398 3072
rect 2410 3068 2411 3072
rect 2413 3068 2414 3072
rect 3239 3068 3240 3072
rect 3242 3068 3245 3072
rect 3247 3068 3248 3072
rect 3260 3068 3261 3072
rect 3263 3068 3264 3072
rect 3276 3068 3277 3072
rect 3279 3068 3282 3072
rect 3284 3068 3285 3072
rect 3302 3068 3303 3072
rect 3305 3068 3306 3072
rect 3318 3068 3319 3072
rect 3321 3068 3322 3072
rect 3334 3068 3335 3072
rect 3337 3068 3340 3072
rect 3342 3068 3343 3072
rect 3355 3068 3356 3072
rect 3358 3068 3359 3072
rect 1511 3038 1512 3042
rect 1514 3038 1517 3042
rect 1519 3038 1520 3042
rect 1532 3038 1533 3042
rect 1535 3038 1536 3042
rect 1548 3038 1549 3042
rect 1551 3038 1554 3042
rect 1556 3038 1557 3042
rect 1574 3038 1575 3042
rect 1577 3038 1578 3042
rect 1590 3038 1591 3042
rect 1593 3038 1594 3042
rect 1606 3038 1607 3042
rect 1609 3038 1612 3042
rect 1614 3038 1615 3042
rect 1627 3038 1628 3042
rect 1630 3038 1631 3042
rect 1643 3038 1644 3042
rect 1646 3038 1649 3042
rect 1651 3038 1652 3042
rect 1664 3038 1665 3042
rect 1667 3038 1668 3042
rect 1680 3038 1681 3042
rect 1683 3038 1686 3042
rect 1688 3038 1689 3042
rect 1706 3038 1707 3042
rect 1709 3038 1710 3042
rect 1722 3038 1723 3042
rect 1725 3038 1726 3042
rect 1738 3038 1739 3042
rect 1741 3038 1744 3042
rect 1746 3038 1747 3042
rect 1759 3038 1760 3042
rect 1762 3038 1763 3042
rect 1775 3038 1776 3042
rect 1778 3038 1781 3042
rect 1783 3038 1784 3042
rect 1796 3038 1797 3042
rect 1799 3038 1800 3042
rect 1812 3038 1813 3042
rect 1815 3038 1818 3042
rect 1820 3038 1821 3042
rect 1838 3038 1839 3042
rect 1841 3038 1842 3042
rect 1854 3038 1855 3042
rect 1857 3038 1858 3042
rect 1870 3038 1871 3042
rect 1873 3038 1876 3042
rect 1878 3038 1879 3042
rect 1891 3038 1892 3042
rect 1894 3038 1895 3042
rect 2456 3038 2457 3042
rect 2459 3038 2462 3042
rect 2464 3038 2465 3042
rect 2477 3038 2478 3042
rect 2480 3038 2481 3042
rect 2493 3038 2494 3042
rect 2496 3038 2499 3042
rect 2501 3038 2502 3042
rect 2519 3038 2520 3042
rect 2522 3038 2523 3042
rect 2535 3038 2536 3042
rect 2538 3038 2539 3042
rect 2551 3038 2552 3042
rect 2554 3038 2557 3042
rect 2559 3038 2560 3042
rect 2572 3038 2573 3042
rect 2575 3038 2576 3042
rect 2588 3038 2589 3042
rect 2591 3038 2594 3042
rect 2596 3038 2597 3042
rect 2609 3038 2610 3042
rect 2612 3038 2613 3042
rect 2625 3038 2626 3042
rect 2628 3038 2631 3042
rect 2633 3038 2634 3042
rect 2651 3038 2652 3042
rect 2654 3038 2655 3042
rect 2667 3038 2668 3042
rect 2670 3038 2671 3042
rect 2683 3038 2684 3042
rect 2686 3038 2689 3042
rect 2691 3038 2692 3042
rect 2704 3038 2705 3042
rect 2707 3038 2708 3042
rect 2720 3038 2721 3042
rect 2723 3038 2726 3042
rect 2728 3038 2729 3042
rect 2741 3038 2742 3042
rect 2744 3038 2745 3042
rect 2757 3038 2758 3042
rect 2760 3038 2763 3042
rect 2765 3038 2766 3042
rect 2783 3038 2784 3042
rect 2786 3038 2787 3042
rect 2799 3038 2800 3042
rect 2802 3038 2803 3042
rect 2815 3038 2816 3042
rect 2818 3038 2821 3042
rect 2823 3038 2824 3042
rect 2836 3038 2837 3042
rect 2839 3038 2840 3042
rect 2436 2994 2440 2995
rect 2436 2991 2440 2992
rect 3381 2994 3385 2995
rect 3381 2991 3385 2992
rect 2294 2982 2295 2986
rect 2297 2982 2300 2986
rect 2302 2982 2303 2986
rect 2315 2982 2316 2986
rect 2318 2982 2319 2986
rect 2331 2982 2332 2986
rect 2334 2982 2337 2986
rect 2339 2982 2340 2986
rect 2357 2982 2358 2986
rect 2360 2982 2361 2986
rect 2373 2982 2374 2986
rect 2376 2982 2377 2986
rect 2389 2982 2390 2986
rect 2392 2982 2395 2986
rect 2397 2982 2398 2986
rect 2410 2982 2411 2986
rect 2413 2982 2414 2986
rect 3239 2982 3240 2986
rect 3242 2982 3245 2986
rect 3247 2982 3248 2986
rect 3260 2982 3261 2986
rect 3263 2982 3264 2986
rect 3276 2982 3277 2986
rect 3279 2982 3282 2986
rect 3284 2982 3285 2986
rect 3302 2982 3303 2986
rect 3305 2982 3306 2986
rect 3318 2982 3319 2986
rect 3321 2982 3322 2986
rect 3334 2982 3335 2986
rect 3337 2982 3340 2986
rect 3342 2982 3343 2986
rect 3355 2982 3356 2986
rect 3358 2982 3359 2986
rect 1511 2952 1512 2956
rect 1514 2952 1517 2956
rect 1519 2952 1520 2956
rect 1532 2952 1533 2956
rect 1535 2952 1536 2956
rect 1548 2952 1549 2956
rect 1551 2952 1554 2956
rect 1556 2952 1557 2956
rect 1574 2952 1575 2956
rect 1577 2952 1578 2956
rect 1590 2952 1591 2956
rect 1593 2952 1594 2956
rect 1606 2952 1607 2956
rect 1609 2952 1612 2956
rect 1614 2952 1615 2956
rect 1627 2952 1628 2956
rect 1630 2952 1631 2956
rect 1643 2952 1644 2956
rect 1646 2952 1649 2956
rect 1651 2952 1652 2956
rect 1664 2952 1665 2956
rect 1667 2952 1668 2956
rect 1680 2952 1681 2956
rect 1683 2952 1686 2956
rect 1688 2952 1689 2956
rect 1706 2952 1707 2956
rect 1709 2952 1710 2956
rect 1722 2952 1723 2956
rect 1725 2952 1726 2956
rect 1738 2952 1739 2956
rect 1741 2952 1744 2956
rect 1746 2952 1747 2956
rect 1759 2952 1760 2956
rect 1762 2952 1763 2956
rect 1775 2952 1776 2956
rect 1778 2952 1781 2956
rect 1783 2952 1784 2956
rect 1796 2952 1797 2956
rect 1799 2952 1800 2956
rect 1812 2952 1813 2956
rect 1815 2952 1818 2956
rect 1820 2952 1821 2956
rect 1838 2952 1839 2956
rect 1841 2952 1842 2956
rect 1854 2952 1855 2956
rect 1857 2952 1858 2956
rect 1870 2952 1871 2956
rect 1873 2952 1876 2956
rect 1878 2952 1879 2956
rect 1891 2952 1892 2956
rect 1894 2952 1895 2956
rect 2456 2952 2457 2956
rect 2459 2952 2462 2956
rect 2464 2952 2465 2956
rect 2477 2952 2478 2956
rect 2480 2952 2481 2956
rect 2493 2952 2494 2956
rect 2496 2952 2499 2956
rect 2501 2952 2502 2956
rect 2519 2952 2520 2956
rect 2522 2952 2523 2956
rect 2535 2952 2536 2956
rect 2538 2952 2539 2956
rect 2551 2952 2552 2956
rect 2554 2952 2557 2956
rect 2559 2952 2560 2956
rect 2572 2952 2573 2956
rect 2575 2952 2576 2956
rect 2588 2952 2589 2956
rect 2591 2952 2594 2956
rect 2596 2952 2597 2956
rect 2609 2952 2610 2956
rect 2612 2952 2613 2956
rect 2625 2952 2626 2956
rect 2628 2952 2631 2956
rect 2633 2952 2634 2956
rect 2651 2952 2652 2956
rect 2654 2952 2655 2956
rect 2667 2952 2668 2956
rect 2670 2952 2671 2956
rect 2683 2952 2684 2956
rect 2686 2952 2689 2956
rect 2691 2952 2692 2956
rect 2704 2952 2705 2956
rect 2707 2952 2708 2956
rect 2720 2952 2721 2956
rect 2723 2952 2726 2956
rect 2728 2952 2729 2956
rect 2741 2952 2742 2956
rect 2744 2952 2745 2956
rect 2757 2952 2758 2956
rect 2760 2952 2763 2956
rect 2765 2952 2766 2956
rect 2783 2952 2784 2956
rect 2786 2952 2787 2956
rect 2799 2952 2800 2956
rect 2802 2952 2803 2956
rect 2815 2952 2816 2956
rect 2818 2952 2821 2956
rect 2823 2952 2824 2956
rect 2836 2952 2837 2956
rect 2839 2952 2840 2956
rect 1743 2908 1744 2912
rect 1746 2908 1747 2912
rect 1767 2908 1768 2912
rect 1770 2908 1771 2912
rect 2688 2908 2689 2912
rect 2691 2908 2692 2912
rect 2712 2908 2713 2912
rect 2715 2908 2716 2912
rect 1763 2897 1764 2901
rect 1766 2897 1767 2901
rect 2708 2897 2709 2901
rect 2711 2897 2712 2901
rect 1755 2885 1759 2886
rect 1755 2882 1759 2883
rect 2700 2885 2704 2886
rect 2700 2882 2704 2883
rect 1743 2874 1744 2878
rect 1746 2874 1747 2878
rect 1767 2874 1768 2878
rect 1770 2874 1771 2878
rect 2688 2874 2689 2878
rect 2691 2874 2692 2878
rect 2712 2874 2713 2878
rect 2715 2874 2716 2878
rect 1511 2812 1512 2816
rect 1514 2812 1517 2816
rect 1519 2812 1520 2816
rect 1532 2812 1533 2816
rect 1535 2812 1536 2816
rect 1548 2812 1549 2816
rect 1551 2812 1554 2816
rect 1556 2812 1557 2816
rect 1574 2812 1575 2816
rect 1577 2812 1578 2816
rect 1590 2812 1591 2816
rect 1593 2812 1594 2816
rect 1606 2812 1607 2816
rect 1609 2812 1612 2816
rect 1614 2812 1615 2816
rect 1627 2812 1628 2816
rect 1630 2812 1631 2816
rect 1643 2812 1644 2816
rect 1646 2812 1649 2816
rect 1651 2812 1652 2816
rect 1664 2812 1665 2816
rect 1667 2812 1668 2816
rect 1680 2812 1681 2816
rect 1683 2812 1686 2816
rect 1688 2812 1689 2816
rect 1706 2812 1707 2816
rect 1709 2812 1710 2816
rect 1722 2812 1723 2816
rect 1725 2812 1726 2816
rect 1738 2812 1739 2816
rect 1741 2812 1744 2816
rect 1746 2812 1747 2816
rect 1759 2812 1760 2816
rect 1762 2812 1763 2816
rect 1775 2812 1776 2816
rect 1778 2812 1781 2816
rect 1783 2812 1784 2816
rect 1796 2812 1797 2816
rect 1799 2812 1800 2816
rect 1812 2812 1813 2816
rect 1815 2812 1818 2816
rect 1820 2812 1821 2816
rect 1838 2812 1839 2816
rect 1841 2812 1842 2816
rect 1854 2812 1855 2816
rect 1857 2812 1858 2816
rect 1870 2812 1871 2816
rect 1873 2812 1876 2816
rect 1878 2812 1879 2816
rect 1891 2812 1892 2816
rect 1894 2812 1895 2816
rect 2456 2812 2457 2816
rect 2459 2812 2462 2816
rect 2464 2812 2465 2816
rect 2477 2812 2478 2816
rect 2480 2812 2481 2816
rect 2493 2812 2494 2816
rect 2496 2812 2499 2816
rect 2501 2812 2502 2816
rect 2519 2812 2520 2816
rect 2522 2812 2523 2816
rect 2535 2812 2536 2816
rect 2538 2812 2539 2816
rect 2551 2812 2552 2816
rect 2554 2812 2557 2816
rect 2559 2812 2560 2816
rect 2572 2812 2573 2816
rect 2575 2812 2576 2816
rect 2588 2812 2589 2816
rect 2591 2812 2594 2816
rect 2596 2812 2597 2816
rect 2609 2812 2610 2816
rect 2612 2812 2613 2816
rect 2625 2812 2626 2816
rect 2628 2812 2631 2816
rect 2633 2812 2634 2816
rect 2651 2812 2652 2816
rect 2654 2812 2655 2816
rect 2667 2812 2668 2816
rect 2670 2812 2671 2816
rect 2683 2812 2684 2816
rect 2686 2812 2689 2816
rect 2691 2812 2692 2816
rect 2704 2812 2705 2816
rect 2707 2812 2708 2816
rect 2720 2812 2721 2816
rect 2723 2812 2726 2816
rect 2728 2812 2729 2816
rect 2741 2812 2742 2816
rect 2744 2812 2745 2816
rect 2757 2812 2758 2816
rect 2760 2812 2763 2816
rect 2765 2812 2766 2816
rect 2783 2812 2784 2816
rect 2786 2812 2787 2816
rect 2799 2812 2800 2816
rect 2802 2812 2803 2816
rect 2815 2812 2816 2816
rect 2818 2812 2821 2816
rect 2823 2812 2824 2816
rect 2836 2812 2837 2816
rect 2839 2812 2840 2816
rect 1995 2733 1996 2737
rect 1998 2733 2001 2737
rect 2003 2733 2004 2737
rect 2016 2733 2017 2737
rect 2019 2733 2020 2737
rect 2032 2733 2033 2737
rect 2035 2733 2038 2737
rect 2040 2733 2041 2737
rect 2058 2733 2059 2737
rect 2061 2733 2062 2737
rect 2074 2733 2075 2737
rect 2077 2733 2078 2737
rect 2090 2733 2091 2737
rect 2093 2733 2096 2737
rect 2098 2733 2099 2737
rect 2111 2733 2112 2737
rect 2114 2733 2115 2737
rect 2127 2733 2128 2737
rect 2130 2733 2133 2737
rect 2135 2733 2136 2737
rect 2148 2733 2149 2737
rect 2151 2733 2152 2737
rect 2164 2733 2165 2737
rect 2167 2733 2170 2737
rect 2172 2733 2173 2737
rect 2190 2733 2191 2737
rect 2193 2733 2194 2737
rect 2206 2733 2207 2737
rect 2209 2733 2210 2737
rect 2222 2733 2223 2737
rect 2225 2733 2228 2737
rect 2230 2733 2231 2737
rect 2243 2733 2244 2737
rect 2246 2733 2247 2737
rect 2259 2733 2260 2737
rect 2262 2733 2265 2737
rect 2267 2733 2268 2737
rect 2280 2733 2281 2737
rect 2283 2733 2284 2737
rect 2296 2733 2297 2737
rect 2299 2733 2302 2737
rect 2304 2733 2305 2737
rect 2322 2733 2323 2737
rect 2325 2733 2326 2737
rect 2338 2733 2339 2737
rect 2341 2733 2342 2737
rect 2354 2733 2355 2737
rect 2357 2733 2360 2737
rect 2362 2733 2363 2737
rect 2375 2733 2376 2737
rect 2378 2733 2379 2737
rect 2391 2733 2392 2737
rect 2394 2733 2397 2737
rect 2399 2733 2400 2737
rect 2412 2733 2413 2737
rect 2415 2733 2416 2737
rect 2428 2733 2429 2737
rect 2431 2733 2434 2737
rect 2436 2733 2437 2737
rect 2454 2733 2455 2737
rect 2457 2733 2458 2737
rect 2470 2733 2471 2737
rect 2473 2733 2474 2737
rect 2486 2733 2487 2737
rect 2489 2733 2492 2737
rect 2494 2733 2495 2737
rect 2507 2733 2508 2737
rect 2510 2733 2511 2737
rect 2940 2733 2941 2737
rect 2943 2733 2946 2737
rect 2948 2733 2949 2737
rect 2961 2733 2962 2737
rect 2964 2733 2965 2737
rect 2977 2733 2978 2737
rect 2980 2733 2983 2737
rect 2985 2733 2986 2737
rect 3003 2733 3004 2737
rect 3006 2733 3007 2737
rect 3019 2733 3020 2737
rect 3022 2733 3023 2737
rect 3035 2733 3036 2737
rect 3038 2733 3041 2737
rect 3043 2733 3044 2737
rect 3056 2733 3057 2737
rect 3059 2733 3060 2737
rect 3072 2733 3073 2737
rect 3075 2733 3078 2737
rect 3080 2733 3081 2737
rect 3093 2733 3094 2737
rect 3096 2733 3097 2737
rect 3109 2733 3110 2737
rect 3112 2733 3115 2737
rect 3117 2733 3118 2737
rect 3135 2733 3136 2737
rect 3138 2733 3139 2737
rect 3151 2733 3152 2737
rect 3154 2733 3155 2737
rect 3167 2733 3168 2737
rect 3170 2733 3173 2737
rect 3175 2733 3176 2737
rect 3188 2733 3189 2737
rect 3191 2733 3192 2737
rect 3204 2733 3205 2737
rect 3207 2733 3210 2737
rect 3212 2733 3213 2737
rect 3225 2733 3226 2737
rect 3228 2733 3229 2737
rect 3241 2733 3242 2737
rect 3244 2733 3247 2737
rect 3249 2733 3250 2737
rect 3267 2733 3268 2737
rect 3270 2733 3271 2737
rect 3283 2733 3284 2737
rect 3286 2733 3287 2737
rect 3299 2733 3300 2737
rect 3302 2733 3305 2737
rect 3307 2733 3308 2737
rect 3320 2733 3321 2737
rect 3323 2733 3324 2737
rect 3336 2733 3337 2737
rect 3339 2733 3342 2737
rect 3344 2733 3345 2737
rect 3357 2733 3358 2737
rect 3360 2733 3361 2737
rect 3373 2733 3374 2737
rect 3376 2733 3379 2737
rect 3381 2733 3382 2737
rect 3399 2733 3400 2737
rect 3402 2733 3403 2737
rect 3415 2733 3416 2737
rect 3418 2733 3419 2737
rect 3431 2733 3432 2737
rect 3434 2733 3437 2737
rect 3439 2733 3440 2737
rect 3452 2733 3453 2737
rect 3455 2733 3456 2737
rect 1643 2700 1644 2704
rect 1646 2700 1649 2704
rect 1651 2700 1652 2704
rect 1664 2700 1665 2704
rect 1667 2700 1668 2704
rect 1680 2700 1681 2704
rect 1683 2700 1686 2704
rect 1688 2700 1689 2704
rect 1706 2700 1707 2704
rect 1709 2700 1710 2704
rect 1722 2700 1723 2704
rect 1725 2700 1726 2704
rect 1738 2700 1739 2704
rect 1741 2700 1744 2704
rect 1746 2700 1747 2704
rect 1759 2700 1760 2704
rect 1762 2700 1763 2704
rect 2588 2700 2589 2704
rect 2591 2700 2594 2704
rect 2596 2700 2597 2704
rect 2609 2700 2610 2704
rect 2612 2700 2613 2704
rect 2625 2700 2626 2704
rect 2628 2700 2631 2704
rect 2633 2700 2634 2704
rect 2651 2700 2652 2704
rect 2654 2700 2655 2704
rect 2667 2700 2668 2704
rect 2670 2700 2671 2704
rect 2683 2700 2684 2704
rect 2686 2700 2689 2704
rect 2691 2700 2692 2704
rect 2704 2700 2705 2704
rect 2707 2700 2708 2704
rect 1767 2663 1768 2667
rect 1770 2663 1771 2667
rect 2174 2667 2175 2671
rect 2177 2667 2178 2671
rect 2198 2663 2201 2667
rect 2203 2663 2206 2667
rect 2208 2663 2209 2667
rect 2255 2667 2256 2671
rect 2258 2667 2259 2671
rect 2279 2663 2282 2667
rect 2284 2663 2287 2667
rect 2289 2663 2290 2667
rect 2228 2659 2229 2663
rect 2231 2659 2232 2663
rect 1650 2654 1651 2658
rect 1653 2654 1654 2658
rect 2000 2654 2001 2658
rect 2003 2654 2004 2658
rect 2016 2654 2017 2658
rect 2019 2654 2020 2658
rect 2032 2654 2033 2658
rect 2035 2654 2036 2658
rect 2051 2654 2056 2658
rect 2058 2654 2061 2658
rect 2063 2654 2064 2658
rect 2085 2654 2087 2658
rect 2089 2654 2090 2658
rect 2107 2654 2108 2658
rect 2110 2654 2111 2658
rect 2123 2654 2128 2658
rect 2130 2654 2133 2658
rect 2135 2654 2136 2658
rect 2150 2654 2151 2658
rect 2153 2654 2154 2658
rect 2309 2659 2310 2663
rect 2312 2659 2313 2663
rect 2712 2663 2713 2667
rect 2715 2663 2716 2667
rect 3119 2667 3120 2671
rect 3122 2667 3123 2671
rect 3143 2663 3146 2667
rect 3148 2663 3151 2667
rect 3153 2663 3154 2667
rect 3200 2667 3201 2671
rect 3203 2667 3204 2671
rect 3224 2663 3227 2667
rect 3229 2663 3232 2667
rect 3234 2663 3235 2667
rect 3173 2659 3174 2663
rect 3176 2659 3177 2663
rect 2595 2654 2596 2658
rect 2598 2654 2599 2658
rect 2945 2654 2946 2658
rect 2948 2654 2949 2658
rect 2961 2654 2962 2658
rect 2964 2654 2965 2658
rect 2977 2654 2978 2658
rect 2980 2654 2981 2658
rect 2996 2654 3001 2658
rect 3003 2654 3006 2658
rect 3008 2654 3009 2658
rect 3030 2654 3032 2658
rect 3034 2654 3035 2658
rect 3052 2654 3053 2658
rect 3055 2654 3056 2658
rect 3068 2654 3073 2658
rect 3075 2654 3078 2658
rect 3080 2654 3081 2658
rect 3095 2654 3096 2658
rect 3098 2654 3099 2658
rect 3254 2659 3255 2663
rect 3257 2659 3258 2663
rect 2000 2608 2001 2612
rect 2003 2608 2004 2612
rect 2016 2608 2017 2612
rect 2019 2608 2020 2612
rect 2032 2608 2033 2612
rect 2035 2608 2036 2612
rect 2051 2608 2056 2612
rect 2058 2608 2061 2612
rect 2063 2608 2064 2612
rect 2085 2608 2087 2612
rect 2089 2608 2090 2612
rect 2107 2608 2108 2612
rect 2110 2608 2111 2612
rect 2123 2608 2128 2612
rect 2130 2608 2133 2612
rect 2135 2608 2136 2612
rect 2150 2608 2151 2612
rect 2153 2608 2154 2612
rect 1634 2598 1635 2602
rect 1637 2598 1638 2602
rect 1650 2598 1651 2602
rect 1653 2598 1656 2602
rect 1658 2598 1659 2602
rect 1671 2598 1672 2602
rect 1674 2598 1675 2602
rect 1687 2598 1688 2602
rect 1690 2598 1691 2602
rect 1708 2598 1709 2602
rect 1711 2598 1714 2602
rect 1716 2598 1717 2602
rect 1729 2598 1730 2602
rect 1732 2598 1733 2602
rect 1745 2598 1746 2602
rect 1748 2598 1751 2602
rect 1753 2598 1754 2602
rect 2198 2607 2201 2611
rect 2203 2607 2206 2611
rect 2208 2607 2209 2611
rect 2279 2607 2282 2611
rect 2284 2607 2287 2611
rect 2289 2607 2290 2611
rect 2945 2608 2946 2612
rect 2948 2608 2949 2612
rect 2961 2608 2962 2612
rect 2964 2608 2965 2612
rect 2977 2608 2978 2612
rect 2980 2608 2981 2612
rect 2996 2608 3001 2612
rect 3003 2608 3006 2612
rect 3008 2608 3009 2612
rect 3030 2608 3032 2612
rect 3034 2608 3035 2612
rect 3052 2608 3053 2612
rect 3055 2608 3056 2612
rect 3068 2608 3073 2612
rect 3075 2608 3078 2612
rect 3080 2608 3081 2612
rect 3095 2608 3096 2612
rect 3098 2608 3099 2612
rect 2579 2598 2580 2602
rect 2582 2598 2583 2602
rect 2595 2598 2596 2602
rect 2598 2598 2601 2602
rect 2603 2598 2604 2602
rect 2616 2598 2617 2602
rect 2619 2598 2620 2602
rect 2632 2598 2633 2602
rect 2635 2598 2636 2602
rect 2653 2598 2654 2602
rect 2656 2598 2659 2602
rect 2661 2598 2662 2602
rect 2674 2598 2675 2602
rect 2677 2598 2678 2602
rect 2690 2598 2691 2602
rect 2693 2598 2696 2602
rect 2698 2598 2699 2602
rect 3143 2607 3146 2611
rect 3148 2607 3151 2611
rect 3153 2607 3154 2611
rect 3224 2607 3227 2611
rect 3229 2607 3232 2611
rect 3234 2607 3235 2611
rect 2198 2531 2201 2535
rect 2203 2531 2206 2535
rect 2208 2531 2209 2535
rect 2279 2535 2280 2539
rect 2282 2535 2283 2539
rect 2303 2531 2306 2535
rect 2308 2531 2311 2535
rect 2313 2531 2314 2535
rect 2228 2527 2229 2531
rect 2231 2527 2232 2531
rect 2000 2522 2001 2526
rect 2003 2522 2004 2526
rect 2016 2522 2017 2526
rect 2019 2522 2020 2526
rect 2032 2522 2033 2526
rect 2035 2522 2036 2526
rect 2051 2522 2056 2526
rect 2058 2522 2061 2526
rect 2063 2522 2064 2526
rect 2085 2522 2087 2526
rect 2089 2522 2090 2526
rect 2107 2522 2108 2526
rect 2110 2522 2111 2526
rect 2123 2522 2128 2526
rect 2130 2522 2133 2526
rect 2135 2522 2136 2526
rect 2150 2522 2151 2526
rect 2153 2522 2154 2526
rect 2333 2527 2334 2531
rect 2336 2527 2337 2531
rect 3143 2531 3146 2535
rect 3148 2531 3151 2535
rect 3153 2531 3154 2535
rect 3224 2535 3225 2539
rect 3227 2535 3228 2539
rect 3248 2531 3251 2535
rect 3253 2531 3256 2535
rect 3258 2531 3259 2535
rect 3173 2527 3174 2531
rect 3176 2527 3177 2531
rect 2945 2522 2946 2526
rect 2948 2522 2949 2526
rect 2961 2522 2962 2526
rect 2964 2522 2965 2526
rect 2977 2522 2978 2526
rect 2980 2522 2981 2526
rect 2996 2522 3001 2526
rect 3003 2522 3006 2526
rect 3008 2522 3009 2526
rect 3030 2522 3032 2526
rect 3034 2522 3035 2526
rect 3052 2522 3053 2526
rect 3055 2522 3056 2526
rect 3068 2522 3073 2526
rect 3075 2522 3078 2526
rect 3080 2522 3081 2526
rect 3095 2522 3096 2526
rect 3098 2522 3099 2526
rect 3278 2527 3279 2531
rect 3281 2527 3282 2531
rect 2000 2476 2001 2480
rect 2003 2476 2004 2480
rect 2016 2476 2017 2480
rect 2019 2476 2020 2480
rect 2032 2476 2033 2480
rect 2035 2476 2036 2480
rect 2051 2476 2056 2480
rect 2058 2476 2061 2480
rect 2063 2476 2064 2480
rect 2085 2476 2087 2480
rect 2089 2476 2090 2480
rect 2107 2476 2108 2480
rect 2110 2476 2111 2480
rect 2123 2476 2128 2480
rect 2130 2476 2133 2480
rect 2135 2476 2136 2480
rect 2150 2476 2151 2480
rect 2153 2476 2154 2480
rect 2198 2476 2201 2480
rect 2203 2476 2206 2480
rect 2208 2476 2209 2480
rect 2303 2476 2306 2480
rect 2308 2476 2311 2480
rect 2313 2476 2314 2480
rect 2945 2476 2946 2480
rect 2948 2476 2949 2480
rect 2961 2476 2962 2480
rect 2964 2476 2965 2480
rect 2977 2476 2978 2480
rect 2980 2476 2981 2480
rect 2996 2476 3001 2480
rect 3003 2476 3006 2480
rect 3008 2476 3009 2480
rect 3030 2476 3032 2480
rect 3034 2476 3035 2480
rect 3052 2476 3053 2480
rect 3055 2476 3056 2480
rect 3068 2476 3073 2480
rect 3075 2476 3078 2480
rect 3080 2476 3081 2480
rect 3095 2476 3096 2480
rect 3098 2476 3099 2480
rect 3143 2476 3146 2480
rect 3148 2476 3151 2480
rect 3153 2476 3154 2480
rect 3248 2476 3251 2480
rect 3253 2476 3256 2480
rect 3258 2476 3259 2480
rect 2198 2399 2201 2403
rect 2203 2399 2206 2403
rect 2208 2399 2209 2403
rect 2255 2403 2256 2407
rect 2258 2403 2259 2407
rect 2279 2399 2282 2403
rect 2284 2399 2287 2403
rect 2289 2399 2290 2403
rect 2345 2403 2346 2407
rect 2348 2403 2349 2407
rect 2369 2399 2372 2403
rect 2374 2399 2377 2403
rect 2379 2399 2380 2403
rect 2228 2395 2229 2399
rect 2231 2395 2232 2399
rect 2000 2390 2001 2394
rect 2003 2390 2004 2394
rect 2016 2390 2017 2394
rect 2019 2390 2020 2394
rect 2032 2390 2033 2394
rect 2035 2390 2036 2394
rect 2051 2390 2056 2394
rect 2058 2390 2061 2394
rect 2063 2390 2064 2394
rect 2085 2390 2087 2394
rect 2089 2390 2090 2394
rect 2107 2390 2108 2394
rect 2110 2390 2111 2394
rect 2123 2390 2128 2394
rect 2130 2390 2133 2394
rect 2135 2390 2136 2394
rect 2150 2390 2151 2394
rect 2153 2390 2154 2394
rect 2309 2395 2310 2399
rect 2312 2395 2313 2399
rect 2399 2395 2400 2399
rect 2402 2395 2403 2399
rect 3143 2399 3146 2403
rect 3148 2399 3151 2403
rect 3153 2399 3154 2403
rect 3200 2403 3201 2407
rect 3203 2403 3204 2407
rect 3224 2399 3227 2403
rect 3229 2399 3232 2403
rect 3234 2399 3235 2403
rect 3290 2403 3291 2407
rect 3293 2403 3294 2407
rect 3314 2399 3317 2403
rect 3319 2399 3322 2403
rect 3324 2399 3325 2403
rect 3173 2395 3174 2399
rect 3176 2395 3177 2399
rect 2945 2390 2946 2394
rect 2948 2390 2949 2394
rect 2961 2390 2962 2394
rect 2964 2390 2965 2394
rect 2977 2390 2978 2394
rect 2980 2390 2981 2394
rect 2996 2390 3001 2394
rect 3003 2390 3006 2394
rect 3008 2390 3009 2394
rect 3030 2390 3032 2394
rect 3034 2390 3035 2394
rect 3052 2390 3053 2394
rect 3055 2390 3056 2394
rect 3068 2390 3073 2394
rect 3075 2390 3078 2394
rect 3080 2390 3081 2394
rect 3095 2390 3096 2394
rect 3098 2390 3099 2394
rect 3254 2395 3255 2399
rect 3257 2395 3258 2399
rect 3344 2395 3345 2399
rect 3347 2395 3348 2399
rect 2000 2344 2001 2348
rect 2003 2344 2004 2348
rect 2016 2344 2017 2348
rect 2019 2344 2020 2348
rect 2032 2344 2033 2348
rect 2035 2344 2036 2348
rect 2051 2344 2056 2348
rect 2058 2344 2061 2348
rect 2063 2344 2064 2348
rect 2085 2344 2087 2348
rect 2089 2344 2090 2348
rect 2107 2344 2108 2348
rect 2110 2344 2111 2348
rect 2123 2344 2128 2348
rect 2130 2344 2133 2348
rect 2135 2344 2136 2348
rect 2150 2344 2151 2348
rect 2153 2344 2154 2348
rect 2198 2341 2201 2345
rect 2203 2341 2206 2345
rect 2208 2341 2209 2345
rect 2279 2341 2282 2345
rect 2284 2341 2287 2345
rect 2289 2341 2290 2345
rect 2369 2341 2372 2345
rect 2374 2341 2377 2345
rect 2379 2341 2380 2345
rect 2945 2344 2946 2348
rect 2948 2344 2949 2348
rect 2961 2344 2962 2348
rect 2964 2344 2965 2348
rect 2977 2344 2978 2348
rect 2980 2344 2981 2348
rect 2996 2344 3001 2348
rect 3003 2344 3006 2348
rect 3008 2344 3009 2348
rect 3030 2344 3032 2348
rect 3034 2344 3035 2348
rect 3052 2344 3053 2348
rect 3055 2344 3056 2348
rect 3068 2344 3073 2348
rect 3075 2344 3078 2348
rect 3080 2344 3081 2348
rect 3095 2344 3096 2348
rect 3098 2344 3099 2348
rect 3143 2341 3146 2345
rect 3148 2341 3151 2345
rect 3153 2341 3154 2345
rect 3224 2341 3227 2345
rect 3229 2341 3232 2345
rect 3234 2341 3235 2345
rect 3314 2341 3317 2345
rect 3319 2341 3322 2345
rect 3324 2341 3325 2345
rect 2198 2267 2201 2271
rect 2203 2267 2206 2271
rect 2208 2267 2209 2271
rect 2228 2263 2229 2267
rect 2231 2263 2232 2267
rect 2000 2258 2001 2262
rect 2003 2258 2004 2262
rect 2016 2258 2017 2262
rect 2019 2258 2020 2262
rect 2032 2258 2033 2262
rect 2035 2258 2036 2262
rect 2051 2258 2056 2262
rect 2058 2258 2061 2262
rect 2063 2258 2064 2262
rect 2085 2258 2087 2262
rect 2089 2258 2090 2262
rect 2107 2258 2108 2262
rect 2110 2258 2111 2262
rect 2123 2258 2128 2262
rect 2130 2258 2133 2262
rect 2135 2258 2136 2262
rect 2150 2258 2151 2262
rect 2153 2258 2154 2262
rect 3143 2267 3146 2271
rect 3148 2267 3151 2271
rect 3153 2267 3154 2271
rect 3173 2263 3174 2267
rect 3176 2263 3177 2267
rect 2945 2258 2946 2262
rect 2948 2258 2949 2262
rect 2961 2258 2962 2262
rect 2964 2258 2965 2262
rect 2977 2258 2978 2262
rect 2980 2258 2981 2262
rect 2996 2258 3001 2262
rect 3003 2258 3006 2262
rect 3008 2258 3009 2262
rect 3030 2258 3032 2262
rect 3034 2258 3035 2262
rect 3052 2258 3053 2262
rect 3055 2258 3056 2262
rect 3068 2258 3073 2262
rect 3075 2258 3078 2262
rect 3080 2258 3081 2262
rect 3095 2258 3096 2262
rect 3098 2258 3099 2262
rect 2000 2212 2001 2216
rect 2003 2212 2004 2216
rect 2016 2212 2017 2216
rect 2019 2212 2020 2216
rect 2032 2212 2033 2216
rect 2035 2212 2036 2216
rect 2051 2212 2056 2216
rect 2058 2212 2061 2216
rect 2063 2212 2064 2216
rect 2085 2212 2087 2216
rect 2089 2212 2090 2216
rect 2107 2212 2108 2216
rect 2110 2212 2111 2216
rect 2123 2212 2128 2216
rect 2130 2212 2133 2216
rect 2135 2212 2136 2216
rect 2150 2212 2151 2216
rect 2153 2212 2154 2216
rect 2234 2212 2235 2216
rect 2237 2212 2238 2216
rect 2242 2212 2248 2216
rect 2252 2212 2253 2216
rect 2255 2212 2256 2216
rect 2277 2212 2278 2216
rect 2280 2212 2281 2216
rect 2293 2212 2294 2216
rect 2296 2212 2297 2216
rect 2312 2212 2317 2216
rect 2319 2212 2322 2216
rect 2324 2212 2325 2216
rect 2346 2212 2348 2216
rect 2350 2212 2351 2216
rect 2368 2212 2369 2216
rect 2371 2212 2372 2216
rect 2384 2212 2389 2216
rect 2391 2212 2394 2216
rect 2396 2212 2397 2216
rect 2411 2212 2412 2216
rect 2414 2212 2415 2216
rect 1511 2198 1512 2202
rect 1514 2198 1517 2202
rect 1519 2198 1520 2202
rect 1532 2198 1533 2202
rect 1535 2198 1536 2202
rect 1548 2198 1549 2202
rect 1551 2198 1554 2202
rect 1556 2198 1557 2202
rect 1574 2198 1575 2202
rect 1577 2198 1578 2202
rect 1590 2198 1591 2202
rect 1593 2198 1594 2202
rect 1606 2198 1607 2202
rect 1609 2198 1612 2202
rect 1614 2198 1615 2202
rect 1627 2198 1628 2202
rect 1630 2198 1631 2202
rect 1643 2198 1644 2202
rect 1646 2198 1649 2202
rect 1651 2198 1652 2202
rect 1664 2198 1665 2202
rect 1667 2198 1668 2202
rect 1680 2198 1681 2202
rect 1683 2198 1686 2202
rect 1688 2198 1689 2202
rect 1706 2198 1707 2202
rect 1709 2198 1710 2202
rect 1722 2198 1723 2202
rect 1725 2198 1726 2202
rect 1738 2198 1739 2202
rect 1741 2198 1744 2202
rect 1746 2198 1747 2202
rect 1759 2198 1760 2202
rect 1762 2198 1763 2202
rect 1775 2198 1776 2202
rect 1778 2198 1781 2202
rect 1783 2198 1784 2202
rect 1796 2198 1797 2202
rect 1799 2198 1800 2202
rect 1812 2198 1813 2202
rect 1815 2198 1818 2202
rect 1820 2198 1821 2202
rect 1838 2198 1839 2202
rect 1841 2198 1842 2202
rect 1854 2198 1855 2202
rect 1857 2198 1858 2202
rect 1870 2198 1871 2202
rect 1873 2198 1876 2202
rect 1878 2198 1879 2202
rect 1891 2198 1892 2202
rect 1894 2198 1895 2202
rect 2198 2205 2201 2209
rect 2203 2205 2206 2209
rect 2208 2205 2209 2209
rect 2945 2212 2946 2216
rect 2948 2212 2949 2216
rect 2961 2212 2962 2216
rect 2964 2212 2965 2216
rect 2977 2212 2978 2216
rect 2980 2212 2981 2216
rect 2996 2212 3001 2216
rect 3003 2212 3006 2216
rect 3008 2212 3009 2216
rect 3030 2212 3032 2216
rect 3034 2212 3035 2216
rect 3052 2212 3053 2216
rect 3055 2212 3056 2216
rect 3068 2212 3073 2216
rect 3075 2212 3078 2216
rect 3080 2212 3081 2216
rect 3095 2212 3096 2216
rect 3098 2212 3099 2216
rect 3179 2212 3180 2216
rect 3182 2212 3183 2216
rect 3187 2212 3193 2216
rect 3197 2212 3198 2216
rect 3200 2212 3201 2216
rect 3222 2212 3223 2216
rect 3225 2212 3226 2216
rect 3238 2212 3239 2216
rect 3241 2212 3242 2216
rect 3257 2212 3262 2216
rect 3264 2212 3267 2216
rect 3269 2212 3270 2216
rect 3291 2212 3293 2216
rect 3295 2212 3296 2216
rect 3313 2212 3314 2216
rect 3316 2212 3317 2216
rect 3329 2212 3334 2216
rect 3336 2212 3339 2216
rect 3341 2212 3342 2216
rect 3356 2212 3357 2216
rect 3359 2212 3360 2216
rect 2456 2198 2457 2202
rect 2459 2198 2462 2202
rect 2464 2198 2465 2202
rect 2477 2198 2478 2202
rect 2480 2198 2481 2202
rect 2493 2198 2494 2202
rect 2496 2198 2499 2202
rect 2501 2198 2502 2202
rect 2519 2198 2520 2202
rect 2522 2198 2523 2202
rect 2535 2198 2536 2202
rect 2538 2198 2539 2202
rect 2551 2198 2552 2202
rect 2554 2198 2557 2202
rect 2559 2198 2560 2202
rect 2572 2198 2573 2202
rect 2575 2198 2576 2202
rect 2588 2198 2589 2202
rect 2591 2198 2594 2202
rect 2596 2198 2597 2202
rect 2609 2198 2610 2202
rect 2612 2198 2613 2202
rect 2625 2198 2626 2202
rect 2628 2198 2631 2202
rect 2633 2198 2634 2202
rect 2651 2198 2652 2202
rect 2654 2198 2655 2202
rect 2667 2198 2668 2202
rect 2670 2198 2671 2202
rect 2683 2198 2684 2202
rect 2686 2198 2689 2202
rect 2691 2198 2692 2202
rect 2704 2198 2705 2202
rect 2707 2198 2708 2202
rect 2720 2198 2721 2202
rect 2723 2198 2726 2202
rect 2728 2198 2729 2202
rect 2741 2198 2742 2202
rect 2744 2198 2745 2202
rect 2757 2198 2758 2202
rect 2760 2198 2763 2202
rect 2765 2198 2766 2202
rect 2783 2198 2784 2202
rect 2786 2198 2787 2202
rect 2799 2198 2800 2202
rect 2802 2198 2803 2202
rect 2815 2198 2816 2202
rect 2818 2198 2821 2202
rect 2823 2198 2824 2202
rect 2836 2198 2837 2202
rect 2839 2198 2840 2202
rect 3143 2205 3146 2209
rect 3148 2205 3151 2209
rect 3153 2205 3154 2209
rect 1626 2154 1627 2158
rect 1629 2154 1630 2158
rect 1650 2154 1651 2158
rect 1653 2154 1654 2158
rect 2424 2158 2428 2159
rect 2424 2155 2428 2156
rect 2571 2154 2572 2158
rect 2574 2154 2575 2158
rect 2595 2154 2596 2158
rect 2598 2154 2599 2158
rect 3369 2158 3373 2159
rect 3369 2155 3373 2156
rect 1646 2141 1647 2145
rect 1649 2141 1650 2145
rect 2591 2141 2592 2145
rect 2594 2141 2595 2145
rect 1638 2129 1642 2130
rect 1638 2126 1642 2127
rect 2583 2129 2587 2130
rect 2583 2126 2587 2127
rect 1626 2118 1627 2122
rect 1629 2118 1630 2122
rect 1650 2118 1651 2122
rect 1653 2118 1654 2122
rect 2571 2118 2572 2122
rect 2574 2118 2575 2122
rect 2595 2118 2596 2122
rect 2598 2118 2599 2122
rect 2294 2086 2295 2090
rect 2297 2086 2300 2090
rect 2302 2086 2303 2090
rect 2315 2086 2316 2090
rect 2318 2086 2319 2090
rect 2331 2086 2332 2090
rect 2334 2086 2337 2090
rect 2339 2086 2340 2090
rect 2357 2086 2358 2090
rect 2360 2086 2361 2090
rect 2373 2086 2374 2090
rect 2376 2086 2377 2090
rect 2389 2086 2390 2090
rect 2392 2086 2395 2090
rect 2397 2086 2398 2090
rect 2410 2086 2411 2090
rect 2413 2086 2414 2090
rect 3239 2086 3240 2090
rect 3242 2086 3245 2090
rect 3247 2086 3248 2090
rect 3260 2086 3261 2090
rect 3263 2086 3264 2090
rect 3276 2086 3277 2090
rect 3279 2086 3282 2090
rect 3284 2086 3285 2090
rect 3302 2086 3303 2090
rect 3305 2086 3306 2090
rect 3318 2086 3319 2090
rect 3321 2086 3322 2090
rect 3334 2086 3335 2090
rect 3337 2086 3340 2090
rect 3342 2086 3343 2090
rect 3355 2086 3356 2090
rect 3358 2086 3359 2090
rect 1511 2056 1512 2060
rect 1514 2056 1517 2060
rect 1519 2056 1520 2060
rect 1532 2056 1533 2060
rect 1535 2056 1536 2060
rect 1548 2056 1549 2060
rect 1551 2056 1554 2060
rect 1556 2056 1557 2060
rect 1574 2056 1575 2060
rect 1577 2056 1578 2060
rect 1590 2056 1591 2060
rect 1593 2056 1594 2060
rect 1606 2056 1607 2060
rect 1609 2056 1612 2060
rect 1614 2056 1615 2060
rect 1627 2056 1628 2060
rect 1630 2056 1631 2060
rect 1643 2056 1644 2060
rect 1646 2056 1649 2060
rect 1651 2056 1652 2060
rect 1664 2056 1665 2060
rect 1667 2056 1668 2060
rect 1680 2056 1681 2060
rect 1683 2056 1686 2060
rect 1688 2056 1689 2060
rect 1706 2056 1707 2060
rect 1709 2056 1710 2060
rect 1722 2056 1723 2060
rect 1725 2056 1726 2060
rect 1738 2056 1739 2060
rect 1741 2056 1744 2060
rect 1746 2056 1747 2060
rect 1759 2056 1760 2060
rect 1762 2056 1763 2060
rect 1775 2056 1776 2060
rect 1778 2056 1781 2060
rect 1783 2056 1784 2060
rect 1796 2056 1797 2060
rect 1799 2056 1800 2060
rect 1812 2056 1813 2060
rect 1815 2056 1818 2060
rect 1820 2056 1821 2060
rect 1838 2056 1839 2060
rect 1841 2056 1842 2060
rect 1854 2056 1855 2060
rect 1857 2056 1858 2060
rect 1870 2056 1871 2060
rect 1873 2056 1876 2060
rect 1878 2056 1879 2060
rect 1891 2056 1892 2060
rect 1894 2056 1895 2060
rect 2456 2056 2457 2060
rect 2459 2056 2462 2060
rect 2464 2056 2465 2060
rect 2477 2056 2478 2060
rect 2480 2056 2481 2060
rect 2493 2056 2494 2060
rect 2496 2056 2499 2060
rect 2501 2056 2502 2060
rect 2519 2056 2520 2060
rect 2522 2056 2523 2060
rect 2535 2056 2536 2060
rect 2538 2056 2539 2060
rect 2551 2056 2552 2060
rect 2554 2056 2557 2060
rect 2559 2056 2560 2060
rect 2572 2056 2573 2060
rect 2575 2056 2576 2060
rect 2588 2056 2589 2060
rect 2591 2056 2594 2060
rect 2596 2056 2597 2060
rect 2609 2056 2610 2060
rect 2612 2056 2613 2060
rect 2625 2056 2626 2060
rect 2628 2056 2631 2060
rect 2633 2056 2634 2060
rect 2651 2056 2652 2060
rect 2654 2056 2655 2060
rect 2667 2056 2668 2060
rect 2670 2056 2671 2060
rect 2683 2056 2684 2060
rect 2686 2056 2689 2060
rect 2691 2056 2692 2060
rect 2704 2056 2705 2060
rect 2707 2056 2708 2060
rect 2720 2056 2721 2060
rect 2723 2056 2726 2060
rect 2728 2056 2729 2060
rect 2741 2056 2742 2060
rect 2744 2056 2745 2060
rect 2757 2056 2758 2060
rect 2760 2056 2763 2060
rect 2765 2056 2766 2060
rect 2783 2056 2784 2060
rect 2786 2056 2787 2060
rect 2799 2056 2800 2060
rect 2802 2056 2803 2060
rect 2815 2056 2816 2060
rect 2818 2056 2821 2060
rect 2823 2056 2824 2060
rect 2836 2056 2837 2060
rect 2839 2056 2840 2060
rect 2436 2012 2440 2013
rect 2436 2009 2440 2010
rect 3381 2012 3385 2013
rect 3381 2009 3385 2010
rect 2294 2000 2295 2004
rect 2297 2000 2300 2004
rect 2302 2000 2303 2004
rect 2315 2000 2316 2004
rect 2318 2000 2319 2004
rect 2331 2000 2332 2004
rect 2334 2000 2337 2004
rect 2339 2000 2340 2004
rect 2357 2000 2358 2004
rect 2360 2000 2361 2004
rect 2373 2000 2374 2004
rect 2376 2000 2377 2004
rect 2389 2000 2390 2004
rect 2392 2000 2395 2004
rect 2397 2000 2398 2004
rect 2410 2000 2411 2004
rect 2413 2000 2414 2004
rect 3239 2000 3240 2004
rect 3242 2000 3245 2004
rect 3247 2000 3248 2004
rect 3260 2000 3261 2004
rect 3263 2000 3264 2004
rect 3276 2000 3277 2004
rect 3279 2000 3282 2004
rect 3284 2000 3285 2004
rect 3302 2000 3303 2004
rect 3305 2000 3306 2004
rect 3318 2000 3319 2004
rect 3321 2000 3322 2004
rect 3334 2000 3335 2004
rect 3337 2000 3340 2004
rect 3342 2000 3343 2004
rect 3355 2000 3356 2004
rect 3358 2000 3359 2004
rect 1511 1970 1512 1974
rect 1514 1970 1517 1974
rect 1519 1970 1520 1974
rect 1532 1970 1533 1974
rect 1535 1970 1536 1974
rect 1548 1970 1549 1974
rect 1551 1970 1554 1974
rect 1556 1970 1557 1974
rect 1574 1970 1575 1974
rect 1577 1970 1578 1974
rect 1590 1970 1591 1974
rect 1593 1970 1594 1974
rect 1606 1970 1607 1974
rect 1609 1970 1612 1974
rect 1614 1970 1615 1974
rect 1627 1970 1628 1974
rect 1630 1970 1631 1974
rect 1643 1970 1644 1974
rect 1646 1970 1649 1974
rect 1651 1970 1652 1974
rect 1664 1970 1665 1974
rect 1667 1970 1668 1974
rect 1680 1970 1681 1974
rect 1683 1970 1686 1974
rect 1688 1970 1689 1974
rect 1706 1970 1707 1974
rect 1709 1970 1710 1974
rect 1722 1970 1723 1974
rect 1725 1970 1726 1974
rect 1738 1970 1739 1974
rect 1741 1970 1744 1974
rect 1746 1970 1747 1974
rect 1759 1970 1760 1974
rect 1762 1970 1763 1974
rect 1775 1970 1776 1974
rect 1778 1970 1781 1974
rect 1783 1970 1784 1974
rect 1796 1970 1797 1974
rect 1799 1970 1800 1974
rect 1812 1970 1813 1974
rect 1815 1970 1818 1974
rect 1820 1970 1821 1974
rect 1838 1970 1839 1974
rect 1841 1970 1842 1974
rect 1854 1970 1855 1974
rect 1857 1970 1858 1974
rect 1870 1970 1871 1974
rect 1873 1970 1876 1974
rect 1878 1970 1879 1974
rect 1891 1970 1892 1974
rect 1894 1970 1895 1974
rect 2456 1970 2457 1974
rect 2459 1970 2462 1974
rect 2464 1970 2465 1974
rect 2477 1970 2478 1974
rect 2480 1970 2481 1974
rect 2493 1970 2494 1974
rect 2496 1970 2499 1974
rect 2501 1970 2502 1974
rect 2519 1970 2520 1974
rect 2522 1970 2523 1974
rect 2535 1970 2536 1974
rect 2538 1970 2539 1974
rect 2551 1970 2552 1974
rect 2554 1970 2557 1974
rect 2559 1970 2560 1974
rect 2572 1970 2573 1974
rect 2575 1970 2576 1974
rect 2588 1970 2589 1974
rect 2591 1970 2594 1974
rect 2596 1970 2597 1974
rect 2609 1970 2610 1974
rect 2612 1970 2613 1974
rect 2625 1970 2626 1974
rect 2628 1970 2631 1974
rect 2633 1970 2634 1974
rect 2651 1970 2652 1974
rect 2654 1970 2655 1974
rect 2667 1970 2668 1974
rect 2670 1970 2671 1974
rect 2683 1970 2684 1974
rect 2686 1970 2689 1974
rect 2691 1970 2692 1974
rect 2704 1970 2705 1974
rect 2707 1970 2708 1974
rect 2720 1970 2721 1974
rect 2723 1970 2726 1974
rect 2728 1970 2729 1974
rect 2741 1970 2742 1974
rect 2744 1970 2745 1974
rect 2757 1970 2758 1974
rect 2760 1970 2763 1974
rect 2765 1970 2766 1974
rect 2783 1970 2784 1974
rect 2786 1970 2787 1974
rect 2799 1970 2800 1974
rect 2802 1970 2803 1974
rect 2815 1970 2816 1974
rect 2818 1970 2821 1974
rect 2823 1970 2824 1974
rect 2836 1970 2837 1974
rect 2839 1970 2840 1974
rect 1743 1926 1744 1930
rect 1746 1926 1747 1930
rect 1767 1926 1768 1930
rect 1770 1926 1771 1930
rect 2688 1926 2689 1930
rect 2691 1926 2692 1930
rect 2712 1926 2713 1930
rect 2715 1926 2716 1930
rect 1763 1915 1764 1919
rect 1766 1915 1767 1919
rect 2708 1915 2709 1919
rect 2711 1915 2712 1919
rect 1755 1903 1759 1904
rect 1755 1900 1759 1901
rect 2700 1903 2704 1904
rect 2700 1900 2704 1901
rect 1743 1892 1744 1896
rect 1746 1892 1747 1896
rect 1767 1892 1768 1896
rect 1770 1892 1771 1896
rect 2688 1892 2689 1896
rect 2691 1892 2692 1896
rect 2712 1892 2713 1896
rect 2715 1892 2716 1896
rect 1511 1830 1512 1834
rect 1514 1830 1517 1834
rect 1519 1830 1520 1834
rect 1532 1830 1533 1834
rect 1535 1830 1536 1834
rect 1548 1830 1549 1834
rect 1551 1830 1554 1834
rect 1556 1830 1557 1834
rect 1574 1830 1575 1834
rect 1577 1830 1578 1834
rect 1590 1830 1591 1834
rect 1593 1830 1594 1834
rect 1606 1830 1607 1834
rect 1609 1830 1612 1834
rect 1614 1830 1615 1834
rect 1627 1830 1628 1834
rect 1630 1830 1631 1834
rect 1643 1830 1644 1834
rect 1646 1830 1649 1834
rect 1651 1830 1652 1834
rect 1664 1830 1665 1834
rect 1667 1830 1668 1834
rect 1680 1830 1681 1834
rect 1683 1830 1686 1834
rect 1688 1830 1689 1834
rect 1706 1830 1707 1834
rect 1709 1830 1710 1834
rect 1722 1830 1723 1834
rect 1725 1830 1726 1834
rect 1738 1830 1739 1834
rect 1741 1830 1744 1834
rect 1746 1830 1747 1834
rect 1759 1830 1760 1834
rect 1762 1830 1763 1834
rect 1775 1830 1776 1834
rect 1778 1830 1781 1834
rect 1783 1830 1784 1834
rect 1796 1830 1797 1834
rect 1799 1830 1800 1834
rect 1812 1830 1813 1834
rect 1815 1830 1818 1834
rect 1820 1830 1821 1834
rect 1838 1830 1839 1834
rect 1841 1830 1842 1834
rect 1854 1830 1855 1834
rect 1857 1830 1858 1834
rect 1870 1830 1871 1834
rect 1873 1830 1876 1834
rect 1878 1830 1879 1834
rect 1891 1830 1892 1834
rect 1894 1830 1895 1834
rect 2456 1830 2457 1834
rect 2459 1830 2462 1834
rect 2464 1830 2465 1834
rect 2477 1830 2478 1834
rect 2480 1830 2481 1834
rect 2493 1830 2494 1834
rect 2496 1830 2499 1834
rect 2501 1830 2502 1834
rect 2519 1830 2520 1834
rect 2522 1830 2523 1834
rect 2535 1830 2536 1834
rect 2538 1830 2539 1834
rect 2551 1830 2552 1834
rect 2554 1830 2557 1834
rect 2559 1830 2560 1834
rect 2572 1830 2573 1834
rect 2575 1830 2576 1834
rect 2588 1830 2589 1834
rect 2591 1830 2594 1834
rect 2596 1830 2597 1834
rect 2609 1830 2610 1834
rect 2612 1830 2613 1834
rect 2625 1830 2626 1834
rect 2628 1830 2631 1834
rect 2633 1830 2634 1834
rect 2651 1830 2652 1834
rect 2654 1830 2655 1834
rect 2667 1830 2668 1834
rect 2670 1830 2671 1834
rect 2683 1830 2684 1834
rect 2686 1830 2689 1834
rect 2691 1830 2692 1834
rect 2704 1830 2705 1834
rect 2707 1830 2708 1834
rect 2720 1830 2721 1834
rect 2723 1830 2726 1834
rect 2728 1830 2729 1834
rect 2741 1830 2742 1834
rect 2744 1830 2745 1834
rect 2757 1830 2758 1834
rect 2760 1830 2763 1834
rect 2765 1830 2766 1834
rect 2783 1830 2784 1834
rect 2786 1830 2787 1834
rect 2799 1830 2800 1834
rect 2802 1830 2803 1834
rect 2815 1830 2816 1834
rect 2818 1830 2821 1834
rect 2823 1830 2824 1834
rect 2836 1830 2837 1834
rect 2839 1830 2840 1834
<< pdiffusion >>
rect 2700 4268 2701 4276
rect 2703 4268 2704 4276
rect 2724 4262 2727 4270
rect 2729 4262 2732 4270
rect 2734 4262 2735 4270
rect 2754 4268 2755 4276
rect 2757 4268 2758 4276
rect 2886 4243 2887 4273
rect 2889 4243 2890 4273
rect 2939 4243 2940 4273
rect 2942 4243 2943 4273
rect 2724 4166 2727 4174
rect 2729 4166 2732 4174
rect 2734 4166 2735 4174
rect 2678 4138 2679 4146
rect 2681 4138 2682 4146
rect 2700 4138 2701 4146
rect 2703 4138 2704 4146
rect 2724 4132 2727 4140
rect 2729 4132 2732 4140
rect 2734 4132 2735 4140
rect 2754 4138 2755 4146
rect 2757 4138 2758 4146
rect 2792 4113 2793 4143
rect 2795 4113 2796 4143
rect 2845 4113 2846 4143
rect 2848 4113 2849 4143
rect 2724 4036 2727 4044
rect 2729 4036 2732 4044
rect 2734 4036 2735 4044
rect 1995 3738 1996 3746
rect 1998 3738 2001 3746
rect 2003 3738 2004 3746
rect 2016 3738 2017 3746
rect 2019 3742 2020 3746
rect 2019 3738 2024 3742
rect 2032 3738 2033 3746
rect 2035 3738 2038 3746
rect 2040 3738 2041 3746
rect 2058 3738 2059 3746
rect 2061 3738 2062 3746
rect 2074 3738 2075 3746
rect 2077 3742 2078 3746
rect 2077 3738 2082 3742
rect 2090 3738 2091 3746
rect 2093 3738 2096 3746
rect 2098 3738 2099 3746
rect 2111 3738 2112 3746
rect 2114 3738 2115 3746
rect 2127 3738 2128 3746
rect 2130 3738 2133 3746
rect 2135 3738 2136 3746
rect 2148 3738 2149 3746
rect 2151 3742 2152 3746
rect 2151 3738 2156 3742
rect 2164 3738 2165 3746
rect 2167 3738 2170 3746
rect 2172 3738 2173 3746
rect 2190 3738 2191 3746
rect 2193 3738 2194 3746
rect 2206 3738 2207 3746
rect 2209 3742 2210 3746
rect 2209 3738 2214 3742
rect 2222 3738 2223 3746
rect 2225 3738 2228 3746
rect 2230 3738 2231 3746
rect 2243 3738 2244 3746
rect 2246 3738 2247 3746
rect 2259 3738 2260 3746
rect 2262 3738 2265 3746
rect 2267 3738 2268 3746
rect 2280 3738 2281 3746
rect 2283 3742 2284 3746
rect 2283 3738 2288 3742
rect 2296 3738 2297 3746
rect 2299 3738 2302 3746
rect 2304 3738 2305 3746
rect 2322 3738 2323 3746
rect 2325 3738 2326 3746
rect 2338 3738 2339 3746
rect 2341 3742 2342 3746
rect 2341 3738 2346 3742
rect 2354 3738 2355 3746
rect 2357 3738 2360 3746
rect 2362 3738 2363 3746
rect 2375 3738 2376 3746
rect 2378 3738 2379 3746
rect 2391 3738 2392 3746
rect 2394 3738 2397 3746
rect 2399 3738 2400 3746
rect 2412 3738 2413 3746
rect 2415 3742 2416 3746
rect 2415 3738 2420 3742
rect 2428 3738 2429 3746
rect 2431 3738 2434 3746
rect 2436 3738 2437 3746
rect 2454 3738 2455 3746
rect 2457 3738 2458 3746
rect 2470 3738 2471 3746
rect 2473 3742 2474 3746
rect 2473 3738 2478 3742
rect 2486 3738 2487 3746
rect 2489 3738 2492 3746
rect 2494 3738 2495 3746
rect 2507 3738 2508 3746
rect 2510 3738 2511 3746
rect 2940 3738 2941 3746
rect 2943 3738 2946 3746
rect 2948 3738 2949 3746
rect 2961 3738 2962 3746
rect 2964 3742 2965 3746
rect 2964 3738 2969 3742
rect 2977 3738 2978 3746
rect 2980 3738 2983 3746
rect 2985 3738 2986 3746
rect 3003 3738 3004 3746
rect 3006 3738 3007 3746
rect 3019 3738 3020 3746
rect 3022 3742 3023 3746
rect 3022 3738 3027 3742
rect 3035 3738 3036 3746
rect 3038 3738 3041 3746
rect 3043 3738 3044 3746
rect 3056 3738 3057 3746
rect 3059 3738 3060 3746
rect 3072 3738 3073 3746
rect 3075 3738 3078 3746
rect 3080 3738 3081 3746
rect 3093 3738 3094 3746
rect 3096 3742 3097 3746
rect 3096 3738 3101 3742
rect 3109 3738 3110 3746
rect 3112 3738 3115 3746
rect 3117 3738 3118 3746
rect 3135 3738 3136 3746
rect 3138 3738 3139 3746
rect 3151 3738 3152 3746
rect 3154 3742 3155 3746
rect 3154 3738 3159 3742
rect 3167 3738 3168 3746
rect 3170 3738 3173 3746
rect 3175 3738 3176 3746
rect 3188 3738 3189 3746
rect 3191 3738 3192 3746
rect 3204 3738 3205 3746
rect 3207 3738 3210 3746
rect 3212 3738 3213 3746
rect 3225 3738 3226 3746
rect 3228 3742 3229 3746
rect 3228 3738 3233 3742
rect 3241 3738 3242 3746
rect 3244 3738 3247 3746
rect 3249 3738 3250 3746
rect 3267 3738 3268 3746
rect 3270 3738 3271 3746
rect 3283 3738 3284 3746
rect 3286 3742 3287 3746
rect 3286 3738 3291 3742
rect 3299 3738 3300 3746
rect 3302 3738 3305 3746
rect 3307 3738 3308 3746
rect 3320 3738 3321 3746
rect 3323 3738 3324 3746
rect 3336 3738 3337 3746
rect 3339 3738 3342 3746
rect 3344 3738 3345 3746
rect 3357 3738 3358 3746
rect 3360 3742 3361 3746
rect 3360 3738 3365 3742
rect 3373 3738 3374 3746
rect 3376 3738 3379 3746
rect 3381 3738 3382 3746
rect 3399 3738 3400 3746
rect 3402 3738 3403 3746
rect 3415 3738 3416 3746
rect 3418 3742 3419 3746
rect 3418 3738 3423 3742
rect 3431 3738 3432 3746
rect 3434 3738 3437 3746
rect 3439 3738 3440 3746
rect 3452 3738 3453 3746
rect 3455 3738 3456 3746
rect 1643 3705 1644 3713
rect 1646 3705 1649 3713
rect 1651 3705 1652 3713
rect 1664 3705 1665 3713
rect 1667 3709 1668 3713
rect 1667 3705 1672 3709
rect 1680 3705 1681 3713
rect 1683 3705 1686 3713
rect 1688 3705 1689 3713
rect 1706 3705 1707 3713
rect 1709 3705 1710 3713
rect 1722 3705 1723 3713
rect 1725 3709 1726 3713
rect 1725 3705 1730 3709
rect 1738 3705 1739 3713
rect 1741 3705 1744 3713
rect 1746 3705 1747 3713
rect 1759 3705 1760 3713
rect 1762 3705 1763 3713
rect 2588 3705 2589 3713
rect 2591 3705 2594 3713
rect 2596 3705 2597 3713
rect 2609 3705 2610 3713
rect 2612 3709 2613 3713
rect 2612 3705 2617 3709
rect 2625 3705 2626 3713
rect 2628 3705 2631 3713
rect 2633 3705 2634 3713
rect 2651 3705 2652 3713
rect 2654 3705 2655 3713
rect 2667 3705 2668 3713
rect 2670 3709 2671 3713
rect 2670 3705 2675 3709
rect 2683 3705 2684 3713
rect 2686 3705 2689 3713
rect 2691 3705 2692 3713
rect 2704 3705 2705 3713
rect 2707 3705 2708 3713
rect 2174 3667 2175 3675
rect 2177 3667 2178 3675
rect 2000 3654 2001 3662
rect 2003 3654 2004 3662
rect 2016 3654 2017 3662
rect 2019 3654 2020 3662
rect 2032 3654 2033 3662
rect 2035 3654 2036 3662
rect 2051 3654 2056 3662
rect 2058 3654 2061 3662
rect 2063 3654 2064 3662
rect 2085 3654 2087 3662
rect 2089 3654 2090 3662
rect 2107 3654 2108 3662
rect 2110 3654 2111 3662
rect 2123 3654 2128 3662
rect 2130 3654 2133 3662
rect 2135 3654 2136 3662
rect 2150 3654 2151 3662
rect 2153 3654 2154 3662
rect 2198 3661 2201 3669
rect 2203 3661 2206 3669
rect 2208 3661 2209 3669
rect 2228 3667 2229 3675
rect 2231 3667 2232 3675
rect 2255 3667 2256 3675
rect 2258 3667 2259 3675
rect 2279 3661 2282 3669
rect 2284 3661 2287 3669
rect 2289 3661 2290 3669
rect 2309 3667 2310 3675
rect 2312 3667 2313 3675
rect 3119 3667 3120 3675
rect 3122 3667 3123 3675
rect 2945 3654 2946 3662
rect 2948 3654 2949 3662
rect 2961 3654 2962 3662
rect 2964 3654 2965 3662
rect 2977 3654 2978 3662
rect 2980 3654 2981 3662
rect 2996 3654 3001 3662
rect 3003 3654 3006 3662
rect 3008 3654 3009 3662
rect 3030 3654 3032 3662
rect 3034 3654 3035 3662
rect 3052 3654 3053 3662
rect 3055 3654 3056 3662
rect 3068 3654 3073 3662
rect 3075 3654 3078 3662
rect 3080 3654 3081 3662
rect 3095 3654 3096 3662
rect 3098 3654 3099 3662
rect 3143 3661 3146 3669
rect 3148 3661 3151 3669
rect 3153 3661 3154 3669
rect 3173 3667 3174 3675
rect 3176 3667 3177 3675
rect 3200 3667 3201 3675
rect 3203 3667 3204 3675
rect 3224 3661 3227 3669
rect 3229 3661 3232 3669
rect 3234 3661 3235 3669
rect 3254 3667 3255 3675
rect 3257 3667 3258 3675
rect 1634 3603 1635 3611
rect 1637 3603 1638 3611
rect 1650 3603 1651 3611
rect 1653 3603 1656 3611
rect 1658 3603 1659 3611
rect 1671 3607 1672 3611
rect 1667 3603 1672 3607
rect 1674 3603 1675 3611
rect 1687 3603 1688 3611
rect 1690 3603 1691 3611
rect 1708 3603 1709 3611
rect 1711 3603 1714 3611
rect 1716 3603 1717 3611
rect 1729 3607 1730 3611
rect 1725 3603 1730 3607
rect 1732 3603 1733 3611
rect 1745 3603 1746 3611
rect 1748 3603 1751 3611
rect 1753 3603 1754 3611
rect 2579 3603 2580 3611
rect 2582 3603 2583 3611
rect 2595 3603 2596 3611
rect 2598 3603 2601 3611
rect 2603 3603 2604 3611
rect 2616 3607 2617 3611
rect 2612 3603 2617 3607
rect 2619 3603 2620 3611
rect 2632 3603 2633 3611
rect 2635 3603 2636 3611
rect 2653 3603 2654 3611
rect 2656 3603 2659 3611
rect 2661 3603 2662 3611
rect 2674 3607 2675 3611
rect 2670 3603 2675 3607
rect 2677 3603 2678 3611
rect 2690 3603 2691 3611
rect 2693 3603 2696 3611
rect 2698 3603 2699 3611
rect 2000 3568 2001 3576
rect 2003 3568 2004 3576
rect 2016 3568 2017 3576
rect 2019 3568 2020 3576
rect 2032 3568 2033 3576
rect 2035 3568 2036 3576
rect 2051 3568 2056 3576
rect 2058 3568 2061 3576
rect 2063 3568 2064 3576
rect 2085 3568 2087 3576
rect 2089 3568 2090 3576
rect 2107 3568 2108 3576
rect 2110 3568 2111 3576
rect 2123 3568 2128 3576
rect 2130 3568 2133 3576
rect 2135 3568 2136 3576
rect 2150 3568 2151 3576
rect 2153 3568 2154 3576
rect 2198 3569 2201 3577
rect 2203 3569 2206 3577
rect 2208 3569 2209 3577
rect 2279 3569 2282 3577
rect 2284 3569 2287 3577
rect 2289 3569 2290 3577
rect 2945 3568 2946 3576
rect 2948 3568 2949 3576
rect 2961 3568 2962 3576
rect 2964 3568 2965 3576
rect 2977 3568 2978 3576
rect 2980 3568 2981 3576
rect 2996 3568 3001 3576
rect 3003 3568 3006 3576
rect 3008 3568 3009 3576
rect 3030 3568 3032 3576
rect 3034 3568 3035 3576
rect 3052 3568 3053 3576
rect 3055 3568 3056 3576
rect 3068 3568 3073 3576
rect 3075 3568 3078 3576
rect 3080 3568 3081 3576
rect 3095 3568 3096 3576
rect 3098 3568 3099 3576
rect 3143 3569 3146 3577
rect 3148 3569 3151 3577
rect 3153 3569 3154 3577
rect 3224 3569 3227 3577
rect 3229 3569 3232 3577
rect 3234 3569 3235 3577
rect 2000 3522 2001 3530
rect 2003 3522 2004 3530
rect 2016 3522 2017 3530
rect 2019 3522 2020 3530
rect 2032 3522 2033 3530
rect 2035 3522 2036 3530
rect 2051 3522 2056 3530
rect 2058 3522 2061 3530
rect 2063 3522 2064 3530
rect 2085 3522 2087 3530
rect 2089 3522 2090 3530
rect 2107 3522 2108 3530
rect 2110 3522 2111 3530
rect 2123 3522 2128 3530
rect 2130 3522 2133 3530
rect 2135 3522 2136 3530
rect 2150 3522 2151 3530
rect 2153 3522 2154 3530
rect 2198 3529 2201 3537
rect 2203 3529 2206 3537
rect 2208 3529 2209 3537
rect 2228 3535 2229 3543
rect 2231 3535 2232 3543
rect 2279 3535 2280 3543
rect 2282 3535 2283 3543
rect 2303 3529 2306 3537
rect 2308 3529 2311 3537
rect 2313 3529 2314 3537
rect 2333 3535 2334 3543
rect 2336 3535 2337 3543
rect 2945 3522 2946 3530
rect 2948 3522 2949 3530
rect 2961 3522 2962 3530
rect 2964 3522 2965 3530
rect 2977 3522 2978 3530
rect 2980 3522 2981 3530
rect 2996 3522 3001 3530
rect 3003 3522 3006 3530
rect 3008 3522 3009 3530
rect 3030 3522 3032 3530
rect 3034 3522 3035 3530
rect 3052 3522 3053 3530
rect 3055 3522 3056 3530
rect 3068 3522 3073 3530
rect 3075 3522 3078 3530
rect 3080 3522 3081 3530
rect 3095 3522 3096 3530
rect 3098 3522 3099 3530
rect 3143 3529 3146 3537
rect 3148 3529 3151 3537
rect 3153 3529 3154 3537
rect 3173 3535 3174 3543
rect 3176 3535 3177 3543
rect 3224 3535 3225 3543
rect 3227 3535 3228 3543
rect 3248 3529 3251 3537
rect 3253 3529 3256 3537
rect 3258 3529 3259 3537
rect 3278 3535 3279 3543
rect 3281 3535 3282 3543
rect 2000 3436 2001 3444
rect 2003 3436 2004 3444
rect 2016 3436 2017 3444
rect 2019 3436 2020 3444
rect 2032 3436 2033 3444
rect 2035 3436 2036 3444
rect 2051 3436 2056 3444
rect 2058 3436 2061 3444
rect 2063 3436 2064 3444
rect 2085 3436 2087 3444
rect 2089 3436 2090 3444
rect 2107 3436 2108 3444
rect 2110 3436 2111 3444
rect 2123 3436 2128 3444
rect 2130 3436 2133 3444
rect 2135 3436 2136 3444
rect 2150 3436 2151 3444
rect 2153 3436 2154 3444
rect 2198 3438 2201 3446
rect 2203 3438 2206 3446
rect 2208 3438 2209 3446
rect 2303 3438 2306 3446
rect 2308 3438 2311 3446
rect 2313 3438 2314 3446
rect 2945 3436 2946 3444
rect 2948 3436 2949 3444
rect 2961 3436 2962 3444
rect 2964 3436 2965 3444
rect 2977 3436 2978 3444
rect 2980 3436 2981 3444
rect 2996 3436 3001 3444
rect 3003 3436 3006 3444
rect 3008 3436 3009 3444
rect 3030 3436 3032 3444
rect 3034 3436 3035 3444
rect 3052 3436 3053 3444
rect 3055 3436 3056 3444
rect 3068 3436 3073 3444
rect 3075 3436 3078 3444
rect 3080 3436 3081 3444
rect 3095 3436 3096 3444
rect 3098 3436 3099 3444
rect 3143 3438 3146 3446
rect 3148 3438 3151 3446
rect 3153 3438 3154 3446
rect 3248 3438 3251 3446
rect 3253 3438 3256 3446
rect 3258 3438 3259 3446
rect 2000 3390 2001 3398
rect 2003 3390 2004 3398
rect 2016 3390 2017 3398
rect 2019 3390 2020 3398
rect 2032 3390 2033 3398
rect 2035 3390 2036 3398
rect 2051 3390 2056 3398
rect 2058 3390 2061 3398
rect 2063 3390 2064 3398
rect 2085 3390 2087 3398
rect 2089 3390 2090 3398
rect 2107 3390 2108 3398
rect 2110 3390 2111 3398
rect 2123 3390 2128 3398
rect 2130 3390 2133 3398
rect 2135 3390 2136 3398
rect 2150 3390 2151 3398
rect 2153 3390 2154 3398
rect 2198 3397 2201 3405
rect 2203 3397 2206 3405
rect 2208 3397 2209 3405
rect 2228 3403 2229 3411
rect 2231 3403 2232 3411
rect 2255 3403 2256 3411
rect 2258 3403 2259 3411
rect 2279 3397 2282 3405
rect 2284 3397 2287 3405
rect 2289 3397 2290 3405
rect 2309 3403 2310 3411
rect 2312 3403 2313 3411
rect 2345 3403 2346 3411
rect 2348 3403 2349 3411
rect 2369 3397 2372 3405
rect 2374 3397 2377 3405
rect 2379 3397 2380 3405
rect 2399 3403 2400 3411
rect 2402 3403 2403 3411
rect 2945 3390 2946 3398
rect 2948 3390 2949 3398
rect 2961 3390 2962 3398
rect 2964 3390 2965 3398
rect 2977 3390 2978 3398
rect 2980 3390 2981 3398
rect 2996 3390 3001 3398
rect 3003 3390 3006 3398
rect 3008 3390 3009 3398
rect 3030 3390 3032 3398
rect 3034 3390 3035 3398
rect 3052 3390 3053 3398
rect 3055 3390 3056 3398
rect 3068 3390 3073 3398
rect 3075 3390 3078 3398
rect 3080 3390 3081 3398
rect 3095 3390 3096 3398
rect 3098 3390 3099 3398
rect 3143 3397 3146 3405
rect 3148 3397 3151 3405
rect 3153 3397 3154 3405
rect 3173 3403 3174 3411
rect 3176 3403 3177 3411
rect 3200 3403 3201 3411
rect 3203 3403 3204 3411
rect 3224 3397 3227 3405
rect 3229 3397 3232 3405
rect 3234 3397 3235 3405
rect 3254 3403 3255 3411
rect 3257 3403 3258 3411
rect 3290 3403 3291 3411
rect 3293 3403 3294 3411
rect 3314 3397 3317 3405
rect 3319 3397 3322 3405
rect 3324 3397 3325 3405
rect 3344 3403 3345 3411
rect 3347 3403 3348 3411
rect 2000 3304 2001 3312
rect 2003 3304 2004 3312
rect 2016 3304 2017 3312
rect 2019 3304 2020 3312
rect 2032 3304 2033 3312
rect 2035 3304 2036 3312
rect 2051 3304 2056 3312
rect 2058 3304 2061 3312
rect 2063 3304 2064 3312
rect 2085 3304 2087 3312
rect 2089 3304 2090 3312
rect 2107 3304 2108 3312
rect 2110 3304 2111 3312
rect 2123 3304 2128 3312
rect 2130 3304 2133 3312
rect 2135 3304 2136 3312
rect 2150 3304 2151 3312
rect 2153 3304 2154 3312
rect 2198 3303 2201 3311
rect 2203 3303 2206 3311
rect 2208 3303 2209 3311
rect 2279 3303 2282 3311
rect 2284 3303 2287 3311
rect 2289 3303 2290 3311
rect 2369 3303 2372 3311
rect 2374 3303 2377 3311
rect 2379 3303 2380 3311
rect 2945 3304 2946 3312
rect 2948 3304 2949 3312
rect 2961 3304 2962 3312
rect 2964 3304 2965 3312
rect 2977 3304 2978 3312
rect 2980 3304 2981 3312
rect 2996 3304 3001 3312
rect 3003 3304 3006 3312
rect 3008 3304 3009 3312
rect 3030 3304 3032 3312
rect 3034 3304 3035 3312
rect 3052 3304 3053 3312
rect 3055 3304 3056 3312
rect 3068 3304 3073 3312
rect 3075 3304 3078 3312
rect 3080 3304 3081 3312
rect 3095 3304 3096 3312
rect 3098 3304 3099 3312
rect 3143 3303 3146 3311
rect 3148 3303 3151 3311
rect 3153 3303 3154 3311
rect 3224 3303 3227 3311
rect 3229 3303 3232 3311
rect 3234 3303 3235 3311
rect 3314 3303 3317 3311
rect 3319 3303 3322 3311
rect 3324 3303 3325 3311
rect 2000 3258 2001 3266
rect 2003 3258 2004 3266
rect 2016 3258 2017 3266
rect 2019 3258 2020 3266
rect 2032 3258 2033 3266
rect 2035 3258 2036 3266
rect 2051 3258 2056 3266
rect 2058 3258 2061 3266
rect 2063 3258 2064 3266
rect 2085 3258 2087 3266
rect 2089 3258 2090 3266
rect 2107 3258 2108 3266
rect 2110 3258 2111 3266
rect 2123 3258 2128 3266
rect 2130 3258 2133 3266
rect 2135 3258 2136 3266
rect 2150 3258 2151 3266
rect 2153 3258 2154 3266
rect 2198 3265 2201 3273
rect 2203 3265 2206 3273
rect 2208 3265 2209 3273
rect 2228 3271 2229 3279
rect 2231 3271 2232 3279
rect 2945 3258 2946 3266
rect 2948 3258 2949 3266
rect 2961 3258 2962 3266
rect 2964 3258 2965 3266
rect 2977 3258 2978 3266
rect 2980 3258 2981 3266
rect 2996 3258 3001 3266
rect 3003 3258 3006 3266
rect 3008 3258 3009 3266
rect 3030 3258 3032 3266
rect 3034 3258 3035 3266
rect 3052 3258 3053 3266
rect 3055 3258 3056 3266
rect 3068 3258 3073 3266
rect 3075 3258 3078 3266
rect 3080 3258 3081 3266
rect 3095 3258 3096 3266
rect 3098 3258 3099 3266
rect 3143 3265 3146 3273
rect 3148 3265 3151 3273
rect 3153 3265 3154 3273
rect 3173 3271 3174 3279
rect 3176 3271 3177 3279
rect 1511 3203 1512 3211
rect 1514 3203 1517 3211
rect 1519 3203 1520 3211
rect 1532 3203 1533 3211
rect 1535 3207 1536 3211
rect 1535 3203 1540 3207
rect 1548 3203 1549 3211
rect 1551 3203 1554 3211
rect 1556 3203 1557 3211
rect 1574 3203 1575 3211
rect 1577 3203 1578 3211
rect 1590 3203 1591 3211
rect 1593 3207 1594 3211
rect 1593 3203 1598 3207
rect 1606 3203 1607 3211
rect 1609 3203 1612 3211
rect 1614 3203 1615 3211
rect 1627 3203 1628 3211
rect 1630 3203 1631 3211
rect 1643 3203 1644 3211
rect 1646 3203 1649 3211
rect 1651 3203 1652 3211
rect 1664 3203 1665 3211
rect 1667 3207 1668 3211
rect 1667 3203 1672 3207
rect 1680 3203 1681 3211
rect 1683 3203 1686 3211
rect 1688 3203 1689 3211
rect 1706 3203 1707 3211
rect 1709 3203 1710 3211
rect 1722 3203 1723 3211
rect 1725 3207 1726 3211
rect 1725 3203 1730 3207
rect 1738 3203 1739 3211
rect 1741 3203 1744 3211
rect 1746 3203 1747 3211
rect 1759 3203 1760 3211
rect 1762 3203 1763 3211
rect 1775 3203 1776 3211
rect 1778 3203 1781 3211
rect 1783 3203 1784 3211
rect 1796 3203 1797 3211
rect 1799 3207 1800 3211
rect 1799 3203 1804 3207
rect 1812 3203 1813 3211
rect 1815 3203 1818 3211
rect 1820 3203 1821 3211
rect 1838 3203 1839 3211
rect 1841 3203 1842 3211
rect 1854 3203 1855 3211
rect 1857 3207 1858 3211
rect 1857 3203 1862 3207
rect 1870 3203 1871 3211
rect 1873 3203 1876 3211
rect 1878 3203 1879 3211
rect 1891 3203 1892 3211
rect 1894 3203 1895 3211
rect 2456 3203 2457 3211
rect 2459 3203 2462 3211
rect 2464 3203 2465 3211
rect 2477 3203 2478 3211
rect 2480 3207 2481 3211
rect 2480 3203 2485 3207
rect 2493 3203 2494 3211
rect 2496 3203 2499 3211
rect 2501 3203 2502 3211
rect 2519 3203 2520 3211
rect 2522 3203 2523 3211
rect 2535 3203 2536 3211
rect 2538 3207 2539 3211
rect 2538 3203 2543 3207
rect 2551 3203 2552 3211
rect 2554 3203 2557 3211
rect 2559 3203 2560 3211
rect 2572 3203 2573 3211
rect 2575 3203 2576 3211
rect 2588 3203 2589 3211
rect 2591 3203 2594 3211
rect 2596 3203 2597 3211
rect 2609 3203 2610 3211
rect 2612 3207 2613 3211
rect 2612 3203 2617 3207
rect 2625 3203 2626 3211
rect 2628 3203 2631 3211
rect 2633 3203 2634 3211
rect 2651 3203 2652 3211
rect 2654 3203 2655 3211
rect 2667 3203 2668 3211
rect 2670 3207 2671 3211
rect 2670 3203 2675 3207
rect 2683 3203 2684 3211
rect 2686 3203 2689 3211
rect 2691 3203 2692 3211
rect 2704 3203 2705 3211
rect 2707 3203 2708 3211
rect 2720 3203 2721 3211
rect 2723 3203 2726 3211
rect 2728 3203 2729 3211
rect 2741 3203 2742 3211
rect 2744 3207 2745 3211
rect 2744 3203 2749 3207
rect 2757 3203 2758 3211
rect 2760 3203 2763 3211
rect 2765 3203 2766 3211
rect 2783 3203 2784 3211
rect 2786 3203 2787 3211
rect 2799 3203 2800 3211
rect 2802 3207 2803 3211
rect 2802 3203 2807 3207
rect 2815 3203 2816 3211
rect 2818 3203 2821 3211
rect 2823 3203 2824 3211
rect 2836 3203 2837 3211
rect 2839 3203 2840 3211
rect 2000 3172 2001 3180
rect 2003 3172 2004 3180
rect 2016 3172 2017 3180
rect 2019 3172 2020 3180
rect 2032 3172 2033 3180
rect 2035 3172 2036 3180
rect 2051 3172 2056 3180
rect 2058 3172 2061 3180
rect 2063 3172 2064 3180
rect 2085 3172 2087 3180
rect 2089 3172 2090 3180
rect 2107 3172 2108 3180
rect 2110 3172 2111 3180
rect 2123 3172 2128 3180
rect 2130 3172 2133 3180
rect 2135 3172 2136 3180
rect 2150 3172 2151 3180
rect 2153 3172 2154 3180
rect 2198 3167 2201 3175
rect 2203 3167 2206 3175
rect 2208 3167 2209 3175
rect 2234 3172 2235 3180
rect 2237 3172 2238 3180
rect 2242 3172 2248 3180
rect 2252 3172 2253 3180
rect 2255 3172 2256 3180
rect 2277 3172 2278 3180
rect 2280 3172 2281 3180
rect 2293 3172 2294 3180
rect 2296 3172 2297 3180
rect 2312 3172 2317 3180
rect 2319 3172 2322 3180
rect 2324 3172 2325 3180
rect 2346 3172 2348 3180
rect 2350 3172 2351 3180
rect 2368 3172 2369 3180
rect 2371 3172 2372 3180
rect 2384 3172 2389 3180
rect 2391 3172 2394 3180
rect 2396 3172 2397 3180
rect 2411 3172 2412 3180
rect 2414 3172 2415 3180
rect 2945 3172 2946 3180
rect 2948 3172 2949 3180
rect 2961 3172 2962 3180
rect 2964 3172 2965 3180
rect 2977 3172 2978 3180
rect 2980 3172 2981 3180
rect 2996 3172 3001 3180
rect 3003 3172 3006 3180
rect 3008 3172 3009 3180
rect 3030 3172 3032 3180
rect 3034 3172 3035 3180
rect 3052 3172 3053 3180
rect 3055 3172 3056 3180
rect 3068 3172 3073 3180
rect 3075 3172 3078 3180
rect 3080 3172 3081 3180
rect 3095 3172 3096 3180
rect 3098 3172 3099 3180
rect 3143 3167 3146 3175
rect 3148 3167 3151 3175
rect 3153 3167 3154 3175
rect 3179 3172 3180 3180
rect 3182 3172 3183 3180
rect 3187 3172 3193 3180
rect 3197 3172 3198 3180
rect 3200 3172 3201 3180
rect 3222 3172 3223 3180
rect 3225 3172 3226 3180
rect 3238 3172 3239 3180
rect 3241 3172 3242 3180
rect 3257 3172 3262 3180
rect 3264 3172 3267 3180
rect 3269 3172 3270 3180
rect 3291 3172 3293 3180
rect 3295 3172 3296 3180
rect 3313 3172 3314 3180
rect 3316 3172 3317 3180
rect 3329 3172 3334 3180
rect 3336 3172 3339 3180
rect 3341 3172 3342 3180
rect 3356 3172 3357 3180
rect 3359 3172 3360 3180
rect 2294 3091 2295 3099
rect 2297 3091 2300 3099
rect 2302 3091 2303 3099
rect 2315 3091 2316 3099
rect 2318 3095 2319 3099
rect 2318 3091 2323 3095
rect 2331 3091 2332 3099
rect 2334 3091 2337 3099
rect 2339 3091 2340 3099
rect 2357 3091 2358 3099
rect 2360 3091 2361 3099
rect 2373 3091 2374 3099
rect 2376 3095 2377 3099
rect 2376 3091 2381 3095
rect 2389 3091 2390 3099
rect 2392 3091 2395 3099
rect 2397 3091 2398 3099
rect 2410 3091 2411 3099
rect 2413 3091 2414 3099
rect 3239 3091 3240 3099
rect 3242 3091 3245 3099
rect 3247 3091 3248 3099
rect 3260 3091 3261 3099
rect 3263 3095 3264 3099
rect 3263 3091 3268 3095
rect 3276 3091 3277 3099
rect 3279 3091 3282 3099
rect 3284 3091 3285 3099
rect 3302 3091 3303 3099
rect 3305 3091 3306 3099
rect 3318 3091 3319 3099
rect 3321 3095 3322 3099
rect 3321 3091 3326 3095
rect 3334 3091 3335 3099
rect 3337 3091 3340 3099
rect 3342 3091 3343 3099
rect 3355 3091 3356 3099
rect 3358 3091 3359 3099
rect 1511 3061 1512 3069
rect 1514 3061 1517 3069
rect 1519 3061 1520 3069
rect 1532 3061 1533 3069
rect 1535 3065 1536 3069
rect 1535 3061 1540 3065
rect 1548 3061 1549 3069
rect 1551 3061 1554 3069
rect 1556 3061 1557 3069
rect 1574 3061 1575 3069
rect 1577 3061 1578 3069
rect 1590 3061 1591 3069
rect 1593 3065 1594 3069
rect 1593 3061 1598 3065
rect 1606 3061 1607 3069
rect 1609 3061 1612 3069
rect 1614 3061 1615 3069
rect 1627 3061 1628 3069
rect 1630 3061 1631 3069
rect 1643 3061 1644 3069
rect 1646 3061 1649 3069
rect 1651 3061 1652 3069
rect 1664 3061 1665 3069
rect 1667 3065 1668 3069
rect 1667 3061 1672 3065
rect 1680 3061 1681 3069
rect 1683 3061 1686 3069
rect 1688 3061 1689 3069
rect 1706 3061 1707 3069
rect 1709 3061 1710 3069
rect 1722 3061 1723 3069
rect 1725 3065 1726 3069
rect 1725 3061 1730 3065
rect 1738 3061 1739 3069
rect 1741 3061 1744 3069
rect 1746 3061 1747 3069
rect 1759 3061 1760 3069
rect 1762 3061 1763 3069
rect 1775 3061 1776 3069
rect 1778 3061 1781 3069
rect 1783 3061 1784 3069
rect 1796 3061 1797 3069
rect 1799 3065 1800 3069
rect 1799 3061 1804 3065
rect 1812 3061 1813 3069
rect 1815 3061 1818 3069
rect 1820 3061 1821 3069
rect 1838 3061 1839 3069
rect 1841 3061 1842 3069
rect 1854 3061 1855 3069
rect 1857 3065 1858 3069
rect 1857 3061 1862 3065
rect 1870 3061 1871 3069
rect 1873 3061 1876 3069
rect 1878 3061 1879 3069
rect 1891 3061 1892 3069
rect 1894 3061 1895 3069
rect 2456 3061 2457 3069
rect 2459 3061 2462 3069
rect 2464 3061 2465 3069
rect 2477 3061 2478 3069
rect 2480 3065 2481 3069
rect 2480 3061 2485 3065
rect 2493 3061 2494 3069
rect 2496 3061 2499 3069
rect 2501 3061 2502 3069
rect 2519 3061 2520 3069
rect 2522 3061 2523 3069
rect 2535 3061 2536 3069
rect 2538 3065 2539 3069
rect 2538 3061 2543 3065
rect 2551 3061 2552 3069
rect 2554 3061 2557 3069
rect 2559 3061 2560 3069
rect 2572 3061 2573 3069
rect 2575 3061 2576 3069
rect 2588 3061 2589 3069
rect 2591 3061 2594 3069
rect 2596 3061 2597 3069
rect 2609 3061 2610 3069
rect 2612 3065 2613 3069
rect 2612 3061 2617 3065
rect 2625 3061 2626 3069
rect 2628 3061 2631 3069
rect 2633 3061 2634 3069
rect 2651 3061 2652 3069
rect 2654 3061 2655 3069
rect 2667 3061 2668 3069
rect 2670 3065 2671 3069
rect 2670 3061 2675 3065
rect 2683 3061 2684 3069
rect 2686 3061 2689 3069
rect 2691 3061 2692 3069
rect 2704 3061 2705 3069
rect 2707 3061 2708 3069
rect 2720 3061 2721 3069
rect 2723 3061 2726 3069
rect 2728 3061 2729 3069
rect 2741 3061 2742 3069
rect 2744 3065 2745 3069
rect 2744 3061 2749 3065
rect 2757 3061 2758 3069
rect 2760 3061 2763 3069
rect 2765 3061 2766 3069
rect 2783 3061 2784 3069
rect 2786 3061 2787 3069
rect 2799 3061 2800 3069
rect 2802 3065 2803 3069
rect 2802 3061 2807 3065
rect 2815 3061 2816 3069
rect 2818 3061 2821 3069
rect 2823 3061 2824 3069
rect 2836 3061 2837 3069
rect 2839 3061 2840 3069
rect 2294 3005 2295 3013
rect 2297 3005 2300 3013
rect 2302 3005 2303 3013
rect 2315 3005 2316 3013
rect 2318 3009 2319 3013
rect 2318 3005 2323 3009
rect 2331 3005 2332 3013
rect 2334 3005 2337 3013
rect 2339 3005 2340 3013
rect 2357 3005 2358 3013
rect 2360 3005 2361 3013
rect 2373 3005 2374 3013
rect 2376 3009 2377 3013
rect 2376 3005 2381 3009
rect 2389 3005 2390 3013
rect 2392 3005 2395 3013
rect 2397 3005 2398 3013
rect 2410 3005 2411 3013
rect 2413 3005 2414 3013
rect 3239 3005 3240 3013
rect 3242 3005 3245 3013
rect 3247 3005 3248 3013
rect 3260 3005 3261 3013
rect 3263 3009 3264 3013
rect 3263 3005 3268 3009
rect 3276 3005 3277 3013
rect 3279 3005 3282 3013
rect 3284 3005 3285 3013
rect 3302 3005 3303 3013
rect 3305 3005 3306 3013
rect 3318 3005 3319 3013
rect 3321 3009 3322 3013
rect 3321 3005 3326 3009
rect 3334 3005 3335 3013
rect 3337 3005 3340 3013
rect 3342 3005 3343 3013
rect 3355 3005 3356 3013
rect 3358 3005 3359 3013
rect 1511 2975 1512 2983
rect 1514 2975 1517 2983
rect 1519 2975 1520 2983
rect 1532 2975 1533 2983
rect 1535 2979 1536 2983
rect 1535 2975 1540 2979
rect 1548 2975 1549 2983
rect 1551 2975 1554 2983
rect 1556 2975 1557 2983
rect 1574 2975 1575 2983
rect 1577 2975 1578 2983
rect 1590 2975 1591 2983
rect 1593 2979 1594 2983
rect 1593 2975 1598 2979
rect 1606 2975 1607 2983
rect 1609 2975 1612 2983
rect 1614 2975 1615 2983
rect 1627 2975 1628 2983
rect 1630 2975 1631 2983
rect 1643 2975 1644 2983
rect 1646 2975 1649 2983
rect 1651 2975 1652 2983
rect 1664 2975 1665 2983
rect 1667 2979 1668 2983
rect 1667 2975 1672 2979
rect 1680 2975 1681 2983
rect 1683 2975 1686 2983
rect 1688 2975 1689 2983
rect 1706 2975 1707 2983
rect 1709 2975 1710 2983
rect 1722 2975 1723 2983
rect 1725 2979 1726 2983
rect 1725 2975 1730 2979
rect 1738 2975 1739 2983
rect 1741 2975 1744 2983
rect 1746 2975 1747 2983
rect 1759 2975 1760 2983
rect 1762 2975 1763 2983
rect 1775 2975 1776 2983
rect 1778 2975 1781 2983
rect 1783 2975 1784 2983
rect 1796 2975 1797 2983
rect 1799 2979 1800 2983
rect 1799 2975 1804 2979
rect 1812 2975 1813 2983
rect 1815 2975 1818 2983
rect 1820 2975 1821 2983
rect 1838 2975 1839 2983
rect 1841 2975 1842 2983
rect 1854 2975 1855 2983
rect 1857 2979 1858 2983
rect 1857 2975 1862 2979
rect 1870 2975 1871 2983
rect 1873 2975 1876 2983
rect 1878 2975 1879 2983
rect 1891 2975 1892 2983
rect 1894 2975 1895 2983
rect 2456 2975 2457 2983
rect 2459 2975 2462 2983
rect 2464 2975 2465 2983
rect 2477 2975 2478 2983
rect 2480 2979 2481 2983
rect 2480 2975 2485 2979
rect 2493 2975 2494 2983
rect 2496 2975 2499 2983
rect 2501 2975 2502 2983
rect 2519 2975 2520 2983
rect 2522 2975 2523 2983
rect 2535 2975 2536 2983
rect 2538 2979 2539 2983
rect 2538 2975 2543 2979
rect 2551 2975 2552 2983
rect 2554 2975 2557 2983
rect 2559 2975 2560 2983
rect 2572 2975 2573 2983
rect 2575 2975 2576 2983
rect 2588 2975 2589 2983
rect 2591 2975 2594 2983
rect 2596 2975 2597 2983
rect 2609 2975 2610 2983
rect 2612 2979 2613 2983
rect 2612 2975 2617 2979
rect 2625 2975 2626 2983
rect 2628 2975 2631 2983
rect 2633 2975 2634 2983
rect 2651 2975 2652 2983
rect 2654 2975 2655 2983
rect 2667 2975 2668 2983
rect 2670 2979 2671 2983
rect 2670 2975 2675 2979
rect 2683 2975 2684 2983
rect 2686 2975 2689 2983
rect 2691 2975 2692 2983
rect 2704 2975 2705 2983
rect 2707 2975 2708 2983
rect 2720 2975 2721 2983
rect 2723 2975 2726 2983
rect 2728 2975 2729 2983
rect 2741 2975 2742 2983
rect 2744 2979 2745 2983
rect 2744 2975 2749 2979
rect 2757 2975 2758 2983
rect 2760 2975 2763 2983
rect 2765 2975 2766 2983
rect 2783 2975 2784 2983
rect 2786 2975 2787 2983
rect 2799 2975 2800 2983
rect 2802 2979 2803 2983
rect 2802 2975 2807 2979
rect 2815 2975 2816 2983
rect 2818 2975 2821 2983
rect 2823 2975 2824 2983
rect 2836 2975 2837 2983
rect 2839 2975 2840 2983
rect 1511 2835 1512 2843
rect 1514 2835 1517 2843
rect 1519 2835 1520 2843
rect 1532 2835 1533 2843
rect 1535 2839 1536 2843
rect 1535 2835 1540 2839
rect 1548 2835 1549 2843
rect 1551 2835 1554 2843
rect 1556 2835 1557 2843
rect 1574 2835 1575 2843
rect 1577 2835 1578 2843
rect 1590 2835 1591 2843
rect 1593 2839 1594 2843
rect 1593 2835 1598 2839
rect 1606 2835 1607 2843
rect 1609 2835 1612 2843
rect 1614 2835 1615 2843
rect 1627 2835 1628 2843
rect 1630 2835 1631 2843
rect 1643 2835 1644 2843
rect 1646 2835 1649 2843
rect 1651 2835 1652 2843
rect 1664 2835 1665 2843
rect 1667 2839 1668 2843
rect 1667 2835 1672 2839
rect 1680 2835 1681 2843
rect 1683 2835 1686 2843
rect 1688 2835 1689 2843
rect 1706 2835 1707 2843
rect 1709 2835 1710 2843
rect 1722 2835 1723 2843
rect 1725 2839 1726 2843
rect 1725 2835 1730 2839
rect 1738 2835 1739 2843
rect 1741 2835 1744 2843
rect 1746 2835 1747 2843
rect 1759 2835 1760 2843
rect 1762 2835 1763 2843
rect 1775 2835 1776 2843
rect 1778 2835 1781 2843
rect 1783 2835 1784 2843
rect 1796 2835 1797 2843
rect 1799 2839 1800 2843
rect 1799 2835 1804 2839
rect 1812 2835 1813 2843
rect 1815 2835 1818 2843
rect 1820 2835 1821 2843
rect 1838 2835 1839 2843
rect 1841 2835 1842 2843
rect 1854 2835 1855 2843
rect 1857 2839 1858 2843
rect 1857 2835 1862 2839
rect 1870 2835 1871 2843
rect 1873 2835 1876 2843
rect 1878 2835 1879 2843
rect 1891 2835 1892 2843
rect 1894 2835 1895 2843
rect 2456 2835 2457 2843
rect 2459 2835 2462 2843
rect 2464 2835 2465 2843
rect 2477 2835 2478 2843
rect 2480 2839 2481 2843
rect 2480 2835 2485 2839
rect 2493 2835 2494 2843
rect 2496 2835 2499 2843
rect 2501 2835 2502 2843
rect 2519 2835 2520 2843
rect 2522 2835 2523 2843
rect 2535 2835 2536 2843
rect 2538 2839 2539 2843
rect 2538 2835 2543 2839
rect 2551 2835 2552 2843
rect 2554 2835 2557 2843
rect 2559 2835 2560 2843
rect 2572 2835 2573 2843
rect 2575 2835 2576 2843
rect 2588 2835 2589 2843
rect 2591 2835 2594 2843
rect 2596 2835 2597 2843
rect 2609 2835 2610 2843
rect 2612 2839 2613 2843
rect 2612 2835 2617 2839
rect 2625 2835 2626 2843
rect 2628 2835 2631 2843
rect 2633 2835 2634 2843
rect 2651 2835 2652 2843
rect 2654 2835 2655 2843
rect 2667 2835 2668 2843
rect 2670 2839 2671 2843
rect 2670 2835 2675 2839
rect 2683 2835 2684 2843
rect 2686 2835 2689 2843
rect 2691 2835 2692 2843
rect 2704 2835 2705 2843
rect 2707 2835 2708 2843
rect 2720 2835 2721 2843
rect 2723 2835 2726 2843
rect 2728 2835 2729 2843
rect 2741 2835 2742 2843
rect 2744 2839 2745 2843
rect 2744 2835 2749 2839
rect 2757 2835 2758 2843
rect 2760 2835 2763 2843
rect 2765 2835 2766 2843
rect 2783 2835 2784 2843
rect 2786 2835 2787 2843
rect 2799 2835 2800 2843
rect 2802 2839 2803 2843
rect 2802 2835 2807 2839
rect 2815 2835 2816 2843
rect 2818 2835 2821 2843
rect 2823 2835 2824 2843
rect 2836 2835 2837 2843
rect 2839 2835 2840 2843
rect 1995 2756 1996 2764
rect 1998 2756 2001 2764
rect 2003 2756 2004 2764
rect 2016 2756 2017 2764
rect 2019 2760 2020 2764
rect 2019 2756 2024 2760
rect 2032 2756 2033 2764
rect 2035 2756 2038 2764
rect 2040 2756 2041 2764
rect 2058 2756 2059 2764
rect 2061 2756 2062 2764
rect 2074 2756 2075 2764
rect 2077 2760 2078 2764
rect 2077 2756 2082 2760
rect 2090 2756 2091 2764
rect 2093 2756 2096 2764
rect 2098 2756 2099 2764
rect 2111 2756 2112 2764
rect 2114 2756 2115 2764
rect 2127 2756 2128 2764
rect 2130 2756 2133 2764
rect 2135 2756 2136 2764
rect 2148 2756 2149 2764
rect 2151 2760 2152 2764
rect 2151 2756 2156 2760
rect 2164 2756 2165 2764
rect 2167 2756 2170 2764
rect 2172 2756 2173 2764
rect 2190 2756 2191 2764
rect 2193 2756 2194 2764
rect 2206 2756 2207 2764
rect 2209 2760 2210 2764
rect 2209 2756 2214 2760
rect 2222 2756 2223 2764
rect 2225 2756 2228 2764
rect 2230 2756 2231 2764
rect 2243 2756 2244 2764
rect 2246 2756 2247 2764
rect 2259 2756 2260 2764
rect 2262 2756 2265 2764
rect 2267 2756 2268 2764
rect 2280 2756 2281 2764
rect 2283 2760 2284 2764
rect 2283 2756 2288 2760
rect 2296 2756 2297 2764
rect 2299 2756 2302 2764
rect 2304 2756 2305 2764
rect 2322 2756 2323 2764
rect 2325 2756 2326 2764
rect 2338 2756 2339 2764
rect 2341 2760 2342 2764
rect 2341 2756 2346 2760
rect 2354 2756 2355 2764
rect 2357 2756 2360 2764
rect 2362 2756 2363 2764
rect 2375 2756 2376 2764
rect 2378 2756 2379 2764
rect 2391 2756 2392 2764
rect 2394 2756 2397 2764
rect 2399 2756 2400 2764
rect 2412 2756 2413 2764
rect 2415 2760 2416 2764
rect 2415 2756 2420 2760
rect 2428 2756 2429 2764
rect 2431 2756 2434 2764
rect 2436 2756 2437 2764
rect 2454 2756 2455 2764
rect 2457 2756 2458 2764
rect 2470 2756 2471 2764
rect 2473 2760 2474 2764
rect 2473 2756 2478 2760
rect 2486 2756 2487 2764
rect 2489 2756 2492 2764
rect 2494 2756 2495 2764
rect 2507 2756 2508 2764
rect 2510 2756 2511 2764
rect 2940 2756 2941 2764
rect 2943 2756 2946 2764
rect 2948 2756 2949 2764
rect 2961 2756 2962 2764
rect 2964 2760 2965 2764
rect 2964 2756 2969 2760
rect 2977 2756 2978 2764
rect 2980 2756 2983 2764
rect 2985 2756 2986 2764
rect 3003 2756 3004 2764
rect 3006 2756 3007 2764
rect 3019 2756 3020 2764
rect 3022 2760 3023 2764
rect 3022 2756 3027 2760
rect 3035 2756 3036 2764
rect 3038 2756 3041 2764
rect 3043 2756 3044 2764
rect 3056 2756 3057 2764
rect 3059 2756 3060 2764
rect 3072 2756 3073 2764
rect 3075 2756 3078 2764
rect 3080 2756 3081 2764
rect 3093 2756 3094 2764
rect 3096 2760 3097 2764
rect 3096 2756 3101 2760
rect 3109 2756 3110 2764
rect 3112 2756 3115 2764
rect 3117 2756 3118 2764
rect 3135 2756 3136 2764
rect 3138 2756 3139 2764
rect 3151 2756 3152 2764
rect 3154 2760 3155 2764
rect 3154 2756 3159 2760
rect 3167 2756 3168 2764
rect 3170 2756 3173 2764
rect 3175 2756 3176 2764
rect 3188 2756 3189 2764
rect 3191 2756 3192 2764
rect 3204 2756 3205 2764
rect 3207 2756 3210 2764
rect 3212 2756 3213 2764
rect 3225 2756 3226 2764
rect 3228 2760 3229 2764
rect 3228 2756 3233 2760
rect 3241 2756 3242 2764
rect 3244 2756 3247 2764
rect 3249 2756 3250 2764
rect 3267 2756 3268 2764
rect 3270 2756 3271 2764
rect 3283 2756 3284 2764
rect 3286 2760 3287 2764
rect 3286 2756 3291 2760
rect 3299 2756 3300 2764
rect 3302 2756 3305 2764
rect 3307 2756 3308 2764
rect 3320 2756 3321 2764
rect 3323 2756 3324 2764
rect 3336 2756 3337 2764
rect 3339 2756 3342 2764
rect 3344 2756 3345 2764
rect 3357 2756 3358 2764
rect 3360 2760 3361 2764
rect 3360 2756 3365 2760
rect 3373 2756 3374 2764
rect 3376 2756 3379 2764
rect 3381 2756 3382 2764
rect 3399 2756 3400 2764
rect 3402 2756 3403 2764
rect 3415 2756 3416 2764
rect 3418 2760 3419 2764
rect 3418 2756 3423 2760
rect 3431 2756 3432 2764
rect 3434 2756 3437 2764
rect 3439 2756 3440 2764
rect 3452 2756 3453 2764
rect 3455 2756 3456 2764
rect 1643 2723 1644 2731
rect 1646 2723 1649 2731
rect 1651 2723 1652 2731
rect 1664 2723 1665 2731
rect 1667 2727 1668 2731
rect 1667 2723 1672 2727
rect 1680 2723 1681 2731
rect 1683 2723 1686 2731
rect 1688 2723 1689 2731
rect 1706 2723 1707 2731
rect 1709 2723 1710 2731
rect 1722 2723 1723 2731
rect 1725 2727 1726 2731
rect 1725 2723 1730 2727
rect 1738 2723 1739 2731
rect 1741 2723 1744 2731
rect 1746 2723 1747 2731
rect 1759 2723 1760 2731
rect 1762 2723 1763 2731
rect 2588 2723 2589 2731
rect 2591 2723 2594 2731
rect 2596 2723 2597 2731
rect 2609 2723 2610 2731
rect 2612 2727 2613 2731
rect 2612 2723 2617 2727
rect 2625 2723 2626 2731
rect 2628 2723 2631 2731
rect 2633 2723 2634 2731
rect 2651 2723 2652 2731
rect 2654 2723 2655 2731
rect 2667 2723 2668 2731
rect 2670 2727 2671 2731
rect 2670 2723 2675 2727
rect 2683 2723 2684 2731
rect 2686 2723 2689 2731
rect 2691 2723 2692 2731
rect 2704 2723 2705 2731
rect 2707 2723 2708 2731
rect 2174 2685 2175 2693
rect 2177 2685 2178 2693
rect 2000 2672 2001 2680
rect 2003 2672 2004 2680
rect 2016 2672 2017 2680
rect 2019 2672 2020 2680
rect 2032 2672 2033 2680
rect 2035 2672 2036 2680
rect 2051 2672 2056 2680
rect 2058 2672 2061 2680
rect 2063 2672 2064 2680
rect 2085 2672 2087 2680
rect 2089 2672 2090 2680
rect 2107 2672 2108 2680
rect 2110 2672 2111 2680
rect 2123 2672 2128 2680
rect 2130 2672 2133 2680
rect 2135 2672 2136 2680
rect 2150 2672 2151 2680
rect 2153 2672 2154 2680
rect 2198 2679 2201 2687
rect 2203 2679 2206 2687
rect 2208 2679 2209 2687
rect 2228 2685 2229 2693
rect 2231 2685 2232 2693
rect 2255 2685 2256 2693
rect 2258 2685 2259 2693
rect 2279 2679 2282 2687
rect 2284 2679 2287 2687
rect 2289 2679 2290 2687
rect 2309 2685 2310 2693
rect 2312 2685 2313 2693
rect 3119 2685 3120 2693
rect 3122 2685 3123 2693
rect 2945 2672 2946 2680
rect 2948 2672 2949 2680
rect 2961 2672 2962 2680
rect 2964 2672 2965 2680
rect 2977 2672 2978 2680
rect 2980 2672 2981 2680
rect 2996 2672 3001 2680
rect 3003 2672 3006 2680
rect 3008 2672 3009 2680
rect 3030 2672 3032 2680
rect 3034 2672 3035 2680
rect 3052 2672 3053 2680
rect 3055 2672 3056 2680
rect 3068 2672 3073 2680
rect 3075 2672 3078 2680
rect 3080 2672 3081 2680
rect 3095 2672 3096 2680
rect 3098 2672 3099 2680
rect 3143 2679 3146 2687
rect 3148 2679 3151 2687
rect 3153 2679 3154 2687
rect 3173 2685 3174 2693
rect 3176 2685 3177 2693
rect 3200 2685 3201 2693
rect 3203 2685 3204 2693
rect 3224 2679 3227 2687
rect 3229 2679 3232 2687
rect 3234 2679 3235 2687
rect 3254 2685 3255 2693
rect 3257 2685 3258 2693
rect 1634 2621 1635 2629
rect 1637 2621 1638 2629
rect 1650 2621 1651 2629
rect 1653 2621 1656 2629
rect 1658 2621 1659 2629
rect 1671 2625 1672 2629
rect 1667 2621 1672 2625
rect 1674 2621 1675 2629
rect 1687 2621 1688 2629
rect 1690 2621 1691 2629
rect 1708 2621 1709 2629
rect 1711 2621 1714 2629
rect 1716 2621 1717 2629
rect 1729 2625 1730 2629
rect 1725 2621 1730 2625
rect 1732 2621 1733 2629
rect 1745 2621 1746 2629
rect 1748 2621 1751 2629
rect 1753 2621 1754 2629
rect 2579 2621 2580 2629
rect 2582 2621 2583 2629
rect 2595 2621 2596 2629
rect 2598 2621 2601 2629
rect 2603 2621 2604 2629
rect 2616 2625 2617 2629
rect 2612 2621 2617 2625
rect 2619 2621 2620 2629
rect 2632 2621 2633 2629
rect 2635 2621 2636 2629
rect 2653 2621 2654 2629
rect 2656 2621 2659 2629
rect 2661 2621 2662 2629
rect 2674 2625 2675 2629
rect 2670 2621 2675 2625
rect 2677 2621 2678 2629
rect 2690 2621 2691 2629
rect 2693 2621 2696 2629
rect 2698 2621 2699 2629
rect 2000 2586 2001 2594
rect 2003 2586 2004 2594
rect 2016 2586 2017 2594
rect 2019 2586 2020 2594
rect 2032 2586 2033 2594
rect 2035 2586 2036 2594
rect 2051 2586 2056 2594
rect 2058 2586 2061 2594
rect 2063 2586 2064 2594
rect 2085 2586 2087 2594
rect 2089 2586 2090 2594
rect 2107 2586 2108 2594
rect 2110 2586 2111 2594
rect 2123 2586 2128 2594
rect 2130 2586 2133 2594
rect 2135 2586 2136 2594
rect 2150 2586 2151 2594
rect 2153 2586 2154 2594
rect 2198 2587 2201 2595
rect 2203 2587 2206 2595
rect 2208 2587 2209 2595
rect 2279 2587 2282 2595
rect 2284 2587 2287 2595
rect 2289 2587 2290 2595
rect 2945 2586 2946 2594
rect 2948 2586 2949 2594
rect 2961 2586 2962 2594
rect 2964 2586 2965 2594
rect 2977 2586 2978 2594
rect 2980 2586 2981 2594
rect 2996 2586 3001 2594
rect 3003 2586 3006 2594
rect 3008 2586 3009 2594
rect 3030 2586 3032 2594
rect 3034 2586 3035 2594
rect 3052 2586 3053 2594
rect 3055 2586 3056 2594
rect 3068 2586 3073 2594
rect 3075 2586 3078 2594
rect 3080 2586 3081 2594
rect 3095 2586 3096 2594
rect 3098 2586 3099 2594
rect 3143 2587 3146 2595
rect 3148 2587 3151 2595
rect 3153 2587 3154 2595
rect 3224 2587 3227 2595
rect 3229 2587 3232 2595
rect 3234 2587 3235 2595
rect 2000 2540 2001 2548
rect 2003 2540 2004 2548
rect 2016 2540 2017 2548
rect 2019 2540 2020 2548
rect 2032 2540 2033 2548
rect 2035 2540 2036 2548
rect 2051 2540 2056 2548
rect 2058 2540 2061 2548
rect 2063 2540 2064 2548
rect 2085 2540 2087 2548
rect 2089 2540 2090 2548
rect 2107 2540 2108 2548
rect 2110 2540 2111 2548
rect 2123 2540 2128 2548
rect 2130 2540 2133 2548
rect 2135 2540 2136 2548
rect 2150 2540 2151 2548
rect 2153 2540 2154 2548
rect 2198 2547 2201 2555
rect 2203 2547 2206 2555
rect 2208 2547 2209 2555
rect 2228 2553 2229 2561
rect 2231 2553 2232 2561
rect 2279 2553 2280 2561
rect 2282 2553 2283 2561
rect 2303 2547 2306 2555
rect 2308 2547 2311 2555
rect 2313 2547 2314 2555
rect 2333 2553 2334 2561
rect 2336 2553 2337 2561
rect 2945 2540 2946 2548
rect 2948 2540 2949 2548
rect 2961 2540 2962 2548
rect 2964 2540 2965 2548
rect 2977 2540 2978 2548
rect 2980 2540 2981 2548
rect 2996 2540 3001 2548
rect 3003 2540 3006 2548
rect 3008 2540 3009 2548
rect 3030 2540 3032 2548
rect 3034 2540 3035 2548
rect 3052 2540 3053 2548
rect 3055 2540 3056 2548
rect 3068 2540 3073 2548
rect 3075 2540 3078 2548
rect 3080 2540 3081 2548
rect 3095 2540 3096 2548
rect 3098 2540 3099 2548
rect 3143 2547 3146 2555
rect 3148 2547 3151 2555
rect 3153 2547 3154 2555
rect 3173 2553 3174 2561
rect 3176 2553 3177 2561
rect 3224 2553 3225 2561
rect 3227 2553 3228 2561
rect 3248 2547 3251 2555
rect 3253 2547 3256 2555
rect 3258 2547 3259 2555
rect 3278 2553 3279 2561
rect 3281 2553 3282 2561
rect 2000 2454 2001 2462
rect 2003 2454 2004 2462
rect 2016 2454 2017 2462
rect 2019 2454 2020 2462
rect 2032 2454 2033 2462
rect 2035 2454 2036 2462
rect 2051 2454 2056 2462
rect 2058 2454 2061 2462
rect 2063 2454 2064 2462
rect 2085 2454 2087 2462
rect 2089 2454 2090 2462
rect 2107 2454 2108 2462
rect 2110 2454 2111 2462
rect 2123 2454 2128 2462
rect 2130 2454 2133 2462
rect 2135 2454 2136 2462
rect 2150 2454 2151 2462
rect 2153 2454 2154 2462
rect 2198 2456 2201 2464
rect 2203 2456 2206 2464
rect 2208 2456 2209 2464
rect 2303 2456 2306 2464
rect 2308 2456 2311 2464
rect 2313 2456 2314 2464
rect 2945 2454 2946 2462
rect 2948 2454 2949 2462
rect 2961 2454 2962 2462
rect 2964 2454 2965 2462
rect 2977 2454 2978 2462
rect 2980 2454 2981 2462
rect 2996 2454 3001 2462
rect 3003 2454 3006 2462
rect 3008 2454 3009 2462
rect 3030 2454 3032 2462
rect 3034 2454 3035 2462
rect 3052 2454 3053 2462
rect 3055 2454 3056 2462
rect 3068 2454 3073 2462
rect 3075 2454 3078 2462
rect 3080 2454 3081 2462
rect 3095 2454 3096 2462
rect 3098 2454 3099 2462
rect 3143 2456 3146 2464
rect 3148 2456 3151 2464
rect 3153 2456 3154 2464
rect 3248 2456 3251 2464
rect 3253 2456 3256 2464
rect 3258 2456 3259 2464
rect 2000 2408 2001 2416
rect 2003 2408 2004 2416
rect 2016 2408 2017 2416
rect 2019 2408 2020 2416
rect 2032 2408 2033 2416
rect 2035 2408 2036 2416
rect 2051 2408 2056 2416
rect 2058 2408 2061 2416
rect 2063 2408 2064 2416
rect 2085 2408 2087 2416
rect 2089 2408 2090 2416
rect 2107 2408 2108 2416
rect 2110 2408 2111 2416
rect 2123 2408 2128 2416
rect 2130 2408 2133 2416
rect 2135 2408 2136 2416
rect 2150 2408 2151 2416
rect 2153 2408 2154 2416
rect 2198 2415 2201 2423
rect 2203 2415 2206 2423
rect 2208 2415 2209 2423
rect 2228 2421 2229 2429
rect 2231 2421 2232 2429
rect 2255 2421 2256 2429
rect 2258 2421 2259 2429
rect 2279 2415 2282 2423
rect 2284 2415 2287 2423
rect 2289 2415 2290 2423
rect 2309 2421 2310 2429
rect 2312 2421 2313 2429
rect 2345 2421 2346 2429
rect 2348 2421 2349 2429
rect 2369 2415 2372 2423
rect 2374 2415 2377 2423
rect 2379 2415 2380 2423
rect 2399 2421 2400 2429
rect 2402 2421 2403 2429
rect 2945 2408 2946 2416
rect 2948 2408 2949 2416
rect 2961 2408 2962 2416
rect 2964 2408 2965 2416
rect 2977 2408 2978 2416
rect 2980 2408 2981 2416
rect 2996 2408 3001 2416
rect 3003 2408 3006 2416
rect 3008 2408 3009 2416
rect 3030 2408 3032 2416
rect 3034 2408 3035 2416
rect 3052 2408 3053 2416
rect 3055 2408 3056 2416
rect 3068 2408 3073 2416
rect 3075 2408 3078 2416
rect 3080 2408 3081 2416
rect 3095 2408 3096 2416
rect 3098 2408 3099 2416
rect 3143 2415 3146 2423
rect 3148 2415 3151 2423
rect 3153 2415 3154 2423
rect 3173 2421 3174 2429
rect 3176 2421 3177 2429
rect 3200 2421 3201 2429
rect 3203 2421 3204 2429
rect 3224 2415 3227 2423
rect 3229 2415 3232 2423
rect 3234 2415 3235 2423
rect 3254 2421 3255 2429
rect 3257 2421 3258 2429
rect 3290 2421 3291 2429
rect 3293 2421 3294 2429
rect 3314 2415 3317 2423
rect 3319 2415 3322 2423
rect 3324 2415 3325 2423
rect 3344 2421 3345 2429
rect 3347 2421 3348 2429
rect 2000 2322 2001 2330
rect 2003 2322 2004 2330
rect 2016 2322 2017 2330
rect 2019 2322 2020 2330
rect 2032 2322 2033 2330
rect 2035 2322 2036 2330
rect 2051 2322 2056 2330
rect 2058 2322 2061 2330
rect 2063 2322 2064 2330
rect 2085 2322 2087 2330
rect 2089 2322 2090 2330
rect 2107 2322 2108 2330
rect 2110 2322 2111 2330
rect 2123 2322 2128 2330
rect 2130 2322 2133 2330
rect 2135 2322 2136 2330
rect 2150 2322 2151 2330
rect 2153 2322 2154 2330
rect 2198 2321 2201 2329
rect 2203 2321 2206 2329
rect 2208 2321 2209 2329
rect 2279 2321 2282 2329
rect 2284 2321 2287 2329
rect 2289 2321 2290 2329
rect 2369 2321 2372 2329
rect 2374 2321 2377 2329
rect 2379 2321 2380 2329
rect 2945 2322 2946 2330
rect 2948 2322 2949 2330
rect 2961 2322 2962 2330
rect 2964 2322 2965 2330
rect 2977 2322 2978 2330
rect 2980 2322 2981 2330
rect 2996 2322 3001 2330
rect 3003 2322 3006 2330
rect 3008 2322 3009 2330
rect 3030 2322 3032 2330
rect 3034 2322 3035 2330
rect 3052 2322 3053 2330
rect 3055 2322 3056 2330
rect 3068 2322 3073 2330
rect 3075 2322 3078 2330
rect 3080 2322 3081 2330
rect 3095 2322 3096 2330
rect 3098 2322 3099 2330
rect 3143 2321 3146 2329
rect 3148 2321 3151 2329
rect 3153 2321 3154 2329
rect 3224 2321 3227 2329
rect 3229 2321 3232 2329
rect 3234 2321 3235 2329
rect 3314 2321 3317 2329
rect 3319 2321 3322 2329
rect 3324 2321 3325 2329
rect 2000 2276 2001 2284
rect 2003 2276 2004 2284
rect 2016 2276 2017 2284
rect 2019 2276 2020 2284
rect 2032 2276 2033 2284
rect 2035 2276 2036 2284
rect 2051 2276 2056 2284
rect 2058 2276 2061 2284
rect 2063 2276 2064 2284
rect 2085 2276 2087 2284
rect 2089 2276 2090 2284
rect 2107 2276 2108 2284
rect 2110 2276 2111 2284
rect 2123 2276 2128 2284
rect 2130 2276 2133 2284
rect 2135 2276 2136 2284
rect 2150 2276 2151 2284
rect 2153 2276 2154 2284
rect 2198 2283 2201 2291
rect 2203 2283 2206 2291
rect 2208 2283 2209 2291
rect 2228 2289 2229 2297
rect 2231 2289 2232 2297
rect 2945 2276 2946 2284
rect 2948 2276 2949 2284
rect 2961 2276 2962 2284
rect 2964 2276 2965 2284
rect 2977 2276 2978 2284
rect 2980 2276 2981 2284
rect 2996 2276 3001 2284
rect 3003 2276 3006 2284
rect 3008 2276 3009 2284
rect 3030 2276 3032 2284
rect 3034 2276 3035 2284
rect 3052 2276 3053 2284
rect 3055 2276 3056 2284
rect 3068 2276 3073 2284
rect 3075 2276 3078 2284
rect 3080 2276 3081 2284
rect 3095 2276 3096 2284
rect 3098 2276 3099 2284
rect 3143 2283 3146 2291
rect 3148 2283 3151 2291
rect 3153 2283 3154 2291
rect 3173 2289 3174 2297
rect 3176 2289 3177 2297
rect 1511 2221 1512 2229
rect 1514 2221 1517 2229
rect 1519 2221 1520 2229
rect 1532 2221 1533 2229
rect 1535 2225 1536 2229
rect 1535 2221 1540 2225
rect 1548 2221 1549 2229
rect 1551 2221 1554 2229
rect 1556 2221 1557 2229
rect 1574 2221 1575 2229
rect 1577 2221 1578 2229
rect 1590 2221 1591 2229
rect 1593 2225 1594 2229
rect 1593 2221 1598 2225
rect 1606 2221 1607 2229
rect 1609 2221 1612 2229
rect 1614 2221 1615 2229
rect 1627 2221 1628 2229
rect 1630 2221 1631 2229
rect 1643 2221 1644 2229
rect 1646 2221 1649 2229
rect 1651 2221 1652 2229
rect 1664 2221 1665 2229
rect 1667 2225 1668 2229
rect 1667 2221 1672 2225
rect 1680 2221 1681 2229
rect 1683 2221 1686 2229
rect 1688 2221 1689 2229
rect 1706 2221 1707 2229
rect 1709 2221 1710 2229
rect 1722 2221 1723 2229
rect 1725 2225 1726 2229
rect 1725 2221 1730 2225
rect 1738 2221 1739 2229
rect 1741 2221 1744 2229
rect 1746 2221 1747 2229
rect 1759 2221 1760 2229
rect 1762 2221 1763 2229
rect 1775 2221 1776 2229
rect 1778 2221 1781 2229
rect 1783 2221 1784 2229
rect 1796 2221 1797 2229
rect 1799 2225 1800 2229
rect 1799 2221 1804 2225
rect 1812 2221 1813 2229
rect 1815 2221 1818 2229
rect 1820 2221 1821 2229
rect 1838 2221 1839 2229
rect 1841 2221 1842 2229
rect 1854 2221 1855 2229
rect 1857 2225 1858 2229
rect 1857 2221 1862 2225
rect 1870 2221 1871 2229
rect 1873 2221 1876 2229
rect 1878 2221 1879 2229
rect 1891 2221 1892 2229
rect 1894 2221 1895 2229
rect 2456 2221 2457 2229
rect 2459 2221 2462 2229
rect 2464 2221 2465 2229
rect 2477 2221 2478 2229
rect 2480 2225 2481 2229
rect 2480 2221 2485 2225
rect 2493 2221 2494 2229
rect 2496 2221 2499 2229
rect 2501 2221 2502 2229
rect 2519 2221 2520 2229
rect 2522 2221 2523 2229
rect 2535 2221 2536 2229
rect 2538 2225 2539 2229
rect 2538 2221 2543 2225
rect 2551 2221 2552 2229
rect 2554 2221 2557 2229
rect 2559 2221 2560 2229
rect 2572 2221 2573 2229
rect 2575 2221 2576 2229
rect 2588 2221 2589 2229
rect 2591 2221 2594 2229
rect 2596 2221 2597 2229
rect 2609 2221 2610 2229
rect 2612 2225 2613 2229
rect 2612 2221 2617 2225
rect 2625 2221 2626 2229
rect 2628 2221 2631 2229
rect 2633 2221 2634 2229
rect 2651 2221 2652 2229
rect 2654 2221 2655 2229
rect 2667 2221 2668 2229
rect 2670 2225 2671 2229
rect 2670 2221 2675 2225
rect 2683 2221 2684 2229
rect 2686 2221 2689 2229
rect 2691 2221 2692 2229
rect 2704 2221 2705 2229
rect 2707 2221 2708 2229
rect 2720 2221 2721 2229
rect 2723 2221 2726 2229
rect 2728 2221 2729 2229
rect 2741 2221 2742 2229
rect 2744 2225 2745 2229
rect 2744 2221 2749 2225
rect 2757 2221 2758 2229
rect 2760 2221 2763 2229
rect 2765 2221 2766 2229
rect 2783 2221 2784 2229
rect 2786 2221 2787 2229
rect 2799 2221 2800 2229
rect 2802 2225 2803 2229
rect 2802 2221 2807 2225
rect 2815 2221 2816 2229
rect 2818 2221 2821 2229
rect 2823 2221 2824 2229
rect 2836 2221 2837 2229
rect 2839 2221 2840 2229
rect 2000 2190 2001 2198
rect 2003 2190 2004 2198
rect 2016 2190 2017 2198
rect 2019 2190 2020 2198
rect 2032 2190 2033 2198
rect 2035 2190 2036 2198
rect 2051 2190 2056 2198
rect 2058 2190 2061 2198
rect 2063 2190 2064 2198
rect 2085 2190 2087 2198
rect 2089 2190 2090 2198
rect 2107 2190 2108 2198
rect 2110 2190 2111 2198
rect 2123 2190 2128 2198
rect 2130 2190 2133 2198
rect 2135 2190 2136 2198
rect 2150 2190 2151 2198
rect 2153 2190 2154 2198
rect 2198 2185 2201 2193
rect 2203 2185 2206 2193
rect 2208 2185 2209 2193
rect 2234 2190 2235 2198
rect 2237 2190 2238 2198
rect 2242 2190 2248 2198
rect 2252 2190 2253 2198
rect 2255 2190 2256 2198
rect 2277 2190 2278 2198
rect 2280 2190 2281 2198
rect 2293 2190 2294 2198
rect 2296 2190 2297 2198
rect 2312 2190 2317 2198
rect 2319 2190 2322 2198
rect 2324 2190 2325 2198
rect 2346 2190 2348 2198
rect 2350 2190 2351 2198
rect 2368 2190 2369 2198
rect 2371 2190 2372 2198
rect 2384 2190 2389 2198
rect 2391 2190 2394 2198
rect 2396 2190 2397 2198
rect 2411 2190 2412 2198
rect 2414 2190 2415 2198
rect 2945 2190 2946 2198
rect 2948 2190 2949 2198
rect 2961 2190 2962 2198
rect 2964 2190 2965 2198
rect 2977 2190 2978 2198
rect 2980 2190 2981 2198
rect 2996 2190 3001 2198
rect 3003 2190 3006 2198
rect 3008 2190 3009 2198
rect 3030 2190 3032 2198
rect 3034 2190 3035 2198
rect 3052 2190 3053 2198
rect 3055 2190 3056 2198
rect 3068 2190 3073 2198
rect 3075 2190 3078 2198
rect 3080 2190 3081 2198
rect 3095 2190 3096 2198
rect 3098 2190 3099 2198
rect 3143 2185 3146 2193
rect 3148 2185 3151 2193
rect 3153 2185 3154 2193
rect 3179 2190 3180 2198
rect 3182 2190 3183 2198
rect 3187 2190 3193 2198
rect 3197 2190 3198 2198
rect 3200 2190 3201 2198
rect 3222 2190 3223 2198
rect 3225 2190 3226 2198
rect 3238 2190 3239 2198
rect 3241 2190 3242 2198
rect 3257 2190 3262 2198
rect 3264 2190 3267 2198
rect 3269 2190 3270 2198
rect 3291 2190 3293 2198
rect 3295 2190 3296 2198
rect 3313 2190 3314 2198
rect 3316 2190 3317 2198
rect 3329 2190 3334 2198
rect 3336 2190 3339 2198
rect 3341 2190 3342 2198
rect 3356 2190 3357 2198
rect 3359 2190 3360 2198
rect 2294 2109 2295 2117
rect 2297 2109 2300 2117
rect 2302 2109 2303 2117
rect 2315 2109 2316 2117
rect 2318 2113 2319 2117
rect 2318 2109 2323 2113
rect 2331 2109 2332 2117
rect 2334 2109 2337 2117
rect 2339 2109 2340 2117
rect 2357 2109 2358 2117
rect 2360 2109 2361 2117
rect 2373 2109 2374 2117
rect 2376 2113 2377 2117
rect 2376 2109 2381 2113
rect 2389 2109 2390 2117
rect 2392 2109 2395 2117
rect 2397 2109 2398 2117
rect 2410 2109 2411 2117
rect 2413 2109 2414 2117
rect 3239 2109 3240 2117
rect 3242 2109 3245 2117
rect 3247 2109 3248 2117
rect 3260 2109 3261 2117
rect 3263 2113 3264 2117
rect 3263 2109 3268 2113
rect 3276 2109 3277 2117
rect 3279 2109 3282 2117
rect 3284 2109 3285 2117
rect 3302 2109 3303 2117
rect 3305 2109 3306 2117
rect 3318 2109 3319 2117
rect 3321 2113 3322 2117
rect 3321 2109 3326 2113
rect 3334 2109 3335 2117
rect 3337 2109 3340 2117
rect 3342 2109 3343 2117
rect 3355 2109 3356 2117
rect 3358 2109 3359 2117
rect 1511 2079 1512 2087
rect 1514 2079 1517 2087
rect 1519 2079 1520 2087
rect 1532 2079 1533 2087
rect 1535 2083 1536 2087
rect 1535 2079 1540 2083
rect 1548 2079 1549 2087
rect 1551 2079 1554 2087
rect 1556 2079 1557 2087
rect 1574 2079 1575 2087
rect 1577 2079 1578 2087
rect 1590 2079 1591 2087
rect 1593 2083 1594 2087
rect 1593 2079 1598 2083
rect 1606 2079 1607 2087
rect 1609 2079 1612 2087
rect 1614 2079 1615 2087
rect 1627 2079 1628 2087
rect 1630 2079 1631 2087
rect 1643 2079 1644 2087
rect 1646 2079 1649 2087
rect 1651 2079 1652 2087
rect 1664 2079 1665 2087
rect 1667 2083 1668 2087
rect 1667 2079 1672 2083
rect 1680 2079 1681 2087
rect 1683 2079 1686 2087
rect 1688 2079 1689 2087
rect 1706 2079 1707 2087
rect 1709 2079 1710 2087
rect 1722 2079 1723 2087
rect 1725 2083 1726 2087
rect 1725 2079 1730 2083
rect 1738 2079 1739 2087
rect 1741 2079 1744 2087
rect 1746 2079 1747 2087
rect 1759 2079 1760 2087
rect 1762 2079 1763 2087
rect 1775 2079 1776 2087
rect 1778 2079 1781 2087
rect 1783 2079 1784 2087
rect 1796 2079 1797 2087
rect 1799 2083 1800 2087
rect 1799 2079 1804 2083
rect 1812 2079 1813 2087
rect 1815 2079 1818 2087
rect 1820 2079 1821 2087
rect 1838 2079 1839 2087
rect 1841 2079 1842 2087
rect 1854 2079 1855 2087
rect 1857 2083 1858 2087
rect 1857 2079 1862 2083
rect 1870 2079 1871 2087
rect 1873 2079 1876 2087
rect 1878 2079 1879 2087
rect 1891 2079 1892 2087
rect 1894 2079 1895 2087
rect 2456 2079 2457 2087
rect 2459 2079 2462 2087
rect 2464 2079 2465 2087
rect 2477 2079 2478 2087
rect 2480 2083 2481 2087
rect 2480 2079 2485 2083
rect 2493 2079 2494 2087
rect 2496 2079 2499 2087
rect 2501 2079 2502 2087
rect 2519 2079 2520 2087
rect 2522 2079 2523 2087
rect 2535 2079 2536 2087
rect 2538 2083 2539 2087
rect 2538 2079 2543 2083
rect 2551 2079 2552 2087
rect 2554 2079 2557 2087
rect 2559 2079 2560 2087
rect 2572 2079 2573 2087
rect 2575 2079 2576 2087
rect 2588 2079 2589 2087
rect 2591 2079 2594 2087
rect 2596 2079 2597 2087
rect 2609 2079 2610 2087
rect 2612 2083 2613 2087
rect 2612 2079 2617 2083
rect 2625 2079 2626 2087
rect 2628 2079 2631 2087
rect 2633 2079 2634 2087
rect 2651 2079 2652 2087
rect 2654 2079 2655 2087
rect 2667 2079 2668 2087
rect 2670 2083 2671 2087
rect 2670 2079 2675 2083
rect 2683 2079 2684 2087
rect 2686 2079 2689 2087
rect 2691 2079 2692 2087
rect 2704 2079 2705 2087
rect 2707 2079 2708 2087
rect 2720 2079 2721 2087
rect 2723 2079 2726 2087
rect 2728 2079 2729 2087
rect 2741 2079 2742 2087
rect 2744 2083 2745 2087
rect 2744 2079 2749 2083
rect 2757 2079 2758 2087
rect 2760 2079 2763 2087
rect 2765 2079 2766 2087
rect 2783 2079 2784 2087
rect 2786 2079 2787 2087
rect 2799 2079 2800 2087
rect 2802 2083 2803 2087
rect 2802 2079 2807 2083
rect 2815 2079 2816 2087
rect 2818 2079 2821 2087
rect 2823 2079 2824 2087
rect 2836 2079 2837 2087
rect 2839 2079 2840 2087
rect 2294 2023 2295 2031
rect 2297 2023 2300 2031
rect 2302 2023 2303 2031
rect 2315 2023 2316 2031
rect 2318 2027 2319 2031
rect 2318 2023 2323 2027
rect 2331 2023 2332 2031
rect 2334 2023 2337 2031
rect 2339 2023 2340 2031
rect 2357 2023 2358 2031
rect 2360 2023 2361 2031
rect 2373 2023 2374 2031
rect 2376 2027 2377 2031
rect 2376 2023 2381 2027
rect 2389 2023 2390 2031
rect 2392 2023 2395 2031
rect 2397 2023 2398 2031
rect 2410 2023 2411 2031
rect 2413 2023 2414 2031
rect 3239 2023 3240 2031
rect 3242 2023 3245 2031
rect 3247 2023 3248 2031
rect 3260 2023 3261 2031
rect 3263 2027 3264 2031
rect 3263 2023 3268 2027
rect 3276 2023 3277 2031
rect 3279 2023 3282 2031
rect 3284 2023 3285 2031
rect 3302 2023 3303 2031
rect 3305 2023 3306 2031
rect 3318 2023 3319 2031
rect 3321 2027 3322 2031
rect 3321 2023 3326 2027
rect 3334 2023 3335 2031
rect 3337 2023 3340 2031
rect 3342 2023 3343 2031
rect 3355 2023 3356 2031
rect 3358 2023 3359 2031
rect 1511 1993 1512 2001
rect 1514 1993 1517 2001
rect 1519 1993 1520 2001
rect 1532 1993 1533 2001
rect 1535 1997 1536 2001
rect 1535 1993 1540 1997
rect 1548 1993 1549 2001
rect 1551 1993 1554 2001
rect 1556 1993 1557 2001
rect 1574 1993 1575 2001
rect 1577 1993 1578 2001
rect 1590 1993 1591 2001
rect 1593 1997 1594 2001
rect 1593 1993 1598 1997
rect 1606 1993 1607 2001
rect 1609 1993 1612 2001
rect 1614 1993 1615 2001
rect 1627 1993 1628 2001
rect 1630 1993 1631 2001
rect 1643 1993 1644 2001
rect 1646 1993 1649 2001
rect 1651 1993 1652 2001
rect 1664 1993 1665 2001
rect 1667 1997 1668 2001
rect 1667 1993 1672 1997
rect 1680 1993 1681 2001
rect 1683 1993 1686 2001
rect 1688 1993 1689 2001
rect 1706 1993 1707 2001
rect 1709 1993 1710 2001
rect 1722 1993 1723 2001
rect 1725 1997 1726 2001
rect 1725 1993 1730 1997
rect 1738 1993 1739 2001
rect 1741 1993 1744 2001
rect 1746 1993 1747 2001
rect 1759 1993 1760 2001
rect 1762 1993 1763 2001
rect 1775 1993 1776 2001
rect 1778 1993 1781 2001
rect 1783 1993 1784 2001
rect 1796 1993 1797 2001
rect 1799 1997 1800 2001
rect 1799 1993 1804 1997
rect 1812 1993 1813 2001
rect 1815 1993 1818 2001
rect 1820 1993 1821 2001
rect 1838 1993 1839 2001
rect 1841 1993 1842 2001
rect 1854 1993 1855 2001
rect 1857 1997 1858 2001
rect 1857 1993 1862 1997
rect 1870 1993 1871 2001
rect 1873 1993 1876 2001
rect 1878 1993 1879 2001
rect 1891 1993 1892 2001
rect 1894 1993 1895 2001
rect 2456 1993 2457 2001
rect 2459 1993 2462 2001
rect 2464 1993 2465 2001
rect 2477 1993 2478 2001
rect 2480 1997 2481 2001
rect 2480 1993 2485 1997
rect 2493 1993 2494 2001
rect 2496 1993 2499 2001
rect 2501 1993 2502 2001
rect 2519 1993 2520 2001
rect 2522 1993 2523 2001
rect 2535 1993 2536 2001
rect 2538 1997 2539 2001
rect 2538 1993 2543 1997
rect 2551 1993 2552 2001
rect 2554 1993 2557 2001
rect 2559 1993 2560 2001
rect 2572 1993 2573 2001
rect 2575 1993 2576 2001
rect 2588 1993 2589 2001
rect 2591 1993 2594 2001
rect 2596 1993 2597 2001
rect 2609 1993 2610 2001
rect 2612 1997 2613 2001
rect 2612 1993 2617 1997
rect 2625 1993 2626 2001
rect 2628 1993 2631 2001
rect 2633 1993 2634 2001
rect 2651 1993 2652 2001
rect 2654 1993 2655 2001
rect 2667 1993 2668 2001
rect 2670 1997 2671 2001
rect 2670 1993 2675 1997
rect 2683 1993 2684 2001
rect 2686 1993 2689 2001
rect 2691 1993 2692 2001
rect 2704 1993 2705 2001
rect 2707 1993 2708 2001
rect 2720 1993 2721 2001
rect 2723 1993 2726 2001
rect 2728 1993 2729 2001
rect 2741 1993 2742 2001
rect 2744 1997 2745 2001
rect 2744 1993 2749 1997
rect 2757 1993 2758 2001
rect 2760 1993 2763 2001
rect 2765 1993 2766 2001
rect 2783 1993 2784 2001
rect 2786 1993 2787 2001
rect 2799 1993 2800 2001
rect 2802 1997 2803 2001
rect 2802 1993 2807 1997
rect 2815 1993 2816 2001
rect 2818 1993 2821 2001
rect 2823 1993 2824 2001
rect 2836 1993 2837 2001
rect 2839 1993 2840 2001
rect 1511 1853 1512 1861
rect 1514 1853 1517 1861
rect 1519 1853 1520 1861
rect 1532 1853 1533 1861
rect 1535 1857 1536 1861
rect 1535 1853 1540 1857
rect 1548 1853 1549 1861
rect 1551 1853 1554 1861
rect 1556 1853 1557 1861
rect 1574 1853 1575 1861
rect 1577 1853 1578 1861
rect 1590 1853 1591 1861
rect 1593 1857 1594 1861
rect 1593 1853 1598 1857
rect 1606 1853 1607 1861
rect 1609 1853 1612 1861
rect 1614 1853 1615 1861
rect 1627 1853 1628 1861
rect 1630 1853 1631 1861
rect 1643 1853 1644 1861
rect 1646 1853 1649 1861
rect 1651 1853 1652 1861
rect 1664 1853 1665 1861
rect 1667 1857 1668 1861
rect 1667 1853 1672 1857
rect 1680 1853 1681 1861
rect 1683 1853 1686 1861
rect 1688 1853 1689 1861
rect 1706 1853 1707 1861
rect 1709 1853 1710 1861
rect 1722 1853 1723 1861
rect 1725 1857 1726 1861
rect 1725 1853 1730 1857
rect 1738 1853 1739 1861
rect 1741 1853 1744 1861
rect 1746 1853 1747 1861
rect 1759 1853 1760 1861
rect 1762 1853 1763 1861
rect 1775 1853 1776 1861
rect 1778 1853 1781 1861
rect 1783 1853 1784 1861
rect 1796 1853 1797 1861
rect 1799 1857 1800 1861
rect 1799 1853 1804 1857
rect 1812 1853 1813 1861
rect 1815 1853 1818 1861
rect 1820 1853 1821 1861
rect 1838 1853 1839 1861
rect 1841 1853 1842 1861
rect 1854 1853 1855 1861
rect 1857 1857 1858 1861
rect 1857 1853 1862 1857
rect 1870 1853 1871 1861
rect 1873 1853 1876 1861
rect 1878 1853 1879 1861
rect 1891 1853 1892 1861
rect 1894 1853 1895 1861
rect 2456 1853 2457 1861
rect 2459 1853 2462 1861
rect 2464 1853 2465 1861
rect 2477 1853 2478 1861
rect 2480 1857 2481 1861
rect 2480 1853 2485 1857
rect 2493 1853 2494 1861
rect 2496 1853 2499 1861
rect 2501 1853 2502 1861
rect 2519 1853 2520 1861
rect 2522 1853 2523 1861
rect 2535 1853 2536 1861
rect 2538 1857 2539 1861
rect 2538 1853 2543 1857
rect 2551 1853 2552 1861
rect 2554 1853 2557 1861
rect 2559 1853 2560 1861
rect 2572 1853 2573 1861
rect 2575 1853 2576 1861
rect 2588 1853 2589 1861
rect 2591 1853 2594 1861
rect 2596 1853 2597 1861
rect 2609 1853 2610 1861
rect 2612 1857 2613 1861
rect 2612 1853 2617 1857
rect 2625 1853 2626 1861
rect 2628 1853 2631 1861
rect 2633 1853 2634 1861
rect 2651 1853 2652 1861
rect 2654 1853 2655 1861
rect 2667 1853 2668 1861
rect 2670 1857 2671 1861
rect 2670 1853 2675 1857
rect 2683 1853 2684 1861
rect 2686 1853 2689 1861
rect 2691 1853 2692 1861
rect 2704 1853 2705 1861
rect 2707 1853 2708 1861
rect 2720 1853 2721 1861
rect 2723 1853 2726 1861
rect 2728 1853 2729 1861
rect 2741 1853 2742 1861
rect 2744 1857 2745 1861
rect 2744 1853 2749 1857
rect 2757 1853 2758 1861
rect 2760 1853 2763 1861
rect 2765 1853 2766 1861
rect 2783 1853 2784 1861
rect 2786 1853 2787 1861
rect 2799 1853 2800 1861
rect 2802 1857 2803 1861
rect 2802 1853 2807 1857
rect 2815 1853 2816 1861
rect 2818 1853 2821 1861
rect 2823 1853 2824 1861
rect 2836 1853 2837 1861
rect 2839 1853 2840 1861
<< ndcontact >>
rect 2696 4250 2700 4254
rect 2704 4250 2708 4254
rect 2720 4246 2724 4250
rect 2735 4246 2739 4250
rect 2750 4242 2754 4246
rect 2758 4242 2762 4246
rect 2870 4211 2886 4223
rect 2890 4211 2906 4223
rect 2923 4211 2939 4223
rect 2943 4211 2959 4223
rect 2720 4186 2724 4190
rect 2735 4186 2739 4190
rect 2674 4120 2678 4124
rect 2682 4120 2686 4124
rect 2696 4120 2700 4124
rect 2704 4120 2708 4124
rect 2720 4116 2724 4120
rect 2735 4116 2739 4120
rect 2750 4112 2754 4116
rect 2758 4112 2762 4116
rect 2776 4081 2792 4093
rect 2796 4081 2812 4093
rect 2829 4081 2845 4093
rect 2849 4081 2865 4093
rect 2720 4056 2724 4060
rect 2735 4056 2739 4060
rect 1991 3715 1995 3719
rect 2004 3715 2008 3719
rect 2012 3715 2016 3719
rect 2020 3715 2024 3719
rect 2028 3715 2032 3719
rect 2041 3715 2045 3719
rect 2054 3715 2058 3719
rect 2062 3715 2066 3719
rect 2070 3715 2074 3719
rect 2078 3715 2082 3719
rect 2086 3715 2090 3719
rect 2099 3715 2103 3719
rect 2107 3715 2111 3719
rect 2115 3715 2119 3719
rect 2123 3715 2127 3719
rect 2136 3715 2140 3719
rect 2144 3715 2148 3719
rect 2152 3715 2156 3719
rect 2160 3715 2164 3719
rect 2173 3715 2177 3719
rect 2186 3715 2190 3719
rect 2194 3715 2198 3719
rect 2202 3715 2206 3719
rect 2210 3715 2214 3719
rect 2218 3715 2222 3719
rect 2231 3715 2235 3719
rect 2239 3715 2243 3719
rect 2247 3715 2251 3719
rect 2255 3715 2259 3719
rect 2268 3715 2272 3719
rect 2276 3715 2280 3719
rect 2284 3715 2288 3719
rect 2292 3715 2296 3719
rect 2305 3715 2309 3719
rect 2318 3715 2322 3719
rect 2326 3715 2330 3719
rect 2334 3715 2338 3719
rect 2342 3715 2346 3719
rect 2350 3715 2354 3719
rect 2363 3715 2367 3719
rect 2371 3715 2375 3719
rect 2379 3715 2383 3719
rect 2387 3715 2391 3719
rect 2400 3715 2404 3719
rect 2408 3715 2412 3719
rect 2416 3715 2420 3719
rect 2424 3715 2428 3719
rect 2437 3715 2441 3719
rect 2450 3715 2454 3719
rect 2458 3715 2462 3719
rect 2466 3715 2470 3719
rect 2474 3715 2478 3719
rect 2482 3715 2486 3719
rect 2495 3715 2499 3719
rect 2503 3715 2507 3719
rect 2511 3715 2515 3719
rect 2936 3715 2940 3719
rect 2949 3715 2953 3719
rect 2957 3715 2961 3719
rect 2965 3715 2969 3719
rect 2973 3715 2977 3719
rect 2986 3715 2990 3719
rect 2999 3715 3003 3719
rect 3007 3715 3011 3719
rect 3015 3715 3019 3719
rect 3023 3715 3027 3719
rect 3031 3715 3035 3719
rect 3044 3715 3048 3719
rect 3052 3715 3056 3719
rect 3060 3715 3064 3719
rect 3068 3715 3072 3719
rect 3081 3715 3085 3719
rect 3089 3715 3093 3719
rect 3097 3715 3101 3719
rect 3105 3715 3109 3719
rect 3118 3715 3122 3719
rect 3131 3715 3135 3719
rect 3139 3715 3143 3719
rect 3147 3715 3151 3719
rect 3155 3715 3159 3719
rect 3163 3715 3167 3719
rect 3176 3715 3180 3719
rect 3184 3715 3188 3719
rect 3192 3715 3196 3719
rect 3200 3715 3204 3719
rect 3213 3715 3217 3719
rect 3221 3715 3225 3719
rect 3229 3715 3233 3719
rect 3237 3715 3241 3719
rect 3250 3715 3254 3719
rect 3263 3715 3267 3719
rect 3271 3715 3275 3719
rect 3279 3715 3283 3719
rect 3287 3715 3291 3719
rect 3295 3715 3299 3719
rect 3308 3715 3312 3719
rect 3316 3715 3320 3719
rect 3324 3715 3328 3719
rect 3332 3715 3336 3719
rect 3345 3715 3349 3719
rect 3353 3715 3357 3719
rect 3361 3715 3365 3719
rect 3369 3715 3373 3719
rect 3382 3715 3386 3719
rect 3395 3715 3399 3719
rect 3403 3715 3407 3719
rect 3411 3715 3415 3719
rect 3419 3715 3423 3719
rect 3427 3715 3431 3719
rect 3440 3715 3444 3719
rect 3448 3715 3452 3719
rect 3456 3715 3460 3719
rect 1639 3682 1643 3686
rect 1652 3682 1656 3686
rect 1660 3682 1664 3686
rect 1668 3682 1672 3686
rect 1676 3682 1680 3686
rect 1689 3682 1693 3686
rect 1702 3682 1706 3686
rect 1710 3682 1714 3686
rect 1718 3682 1722 3686
rect 1726 3682 1730 3686
rect 1734 3682 1738 3686
rect 1747 3682 1751 3686
rect 1755 3682 1759 3686
rect 1763 3682 1767 3686
rect 2584 3682 2588 3686
rect 2597 3682 2601 3686
rect 2605 3682 2609 3686
rect 2613 3682 2617 3686
rect 2621 3682 2625 3686
rect 2634 3682 2638 3686
rect 2647 3682 2651 3686
rect 2655 3682 2659 3686
rect 2663 3682 2667 3686
rect 2671 3682 2675 3686
rect 2679 3682 2683 3686
rect 2692 3682 2696 3686
rect 2700 3682 2704 3686
rect 2708 3682 2712 3686
rect 1763 3645 1767 3649
rect 1771 3645 1775 3649
rect 2170 3649 2174 3653
rect 2178 3649 2182 3653
rect 2194 3645 2198 3649
rect 2209 3645 2213 3649
rect 2251 3649 2255 3653
rect 2259 3649 2263 3653
rect 2275 3645 2279 3649
rect 2290 3645 2294 3649
rect 2224 3641 2228 3645
rect 2232 3641 2236 3645
rect 1646 3636 1650 3640
rect 1654 3636 1658 3640
rect 1996 3636 2000 3640
rect 2004 3636 2008 3640
rect 2012 3636 2016 3640
rect 2020 3636 2024 3640
rect 2028 3636 2032 3640
rect 2036 3636 2040 3640
rect 2047 3636 2051 3640
rect 2064 3636 2068 3640
rect 2081 3636 2085 3640
rect 2090 3636 2094 3640
rect 2103 3636 2107 3640
rect 2111 3636 2115 3640
rect 2119 3636 2123 3640
rect 2136 3636 2140 3640
rect 2146 3636 2150 3640
rect 2154 3636 2158 3640
rect 2305 3641 2309 3645
rect 2313 3641 2317 3645
rect 2708 3645 2712 3649
rect 2716 3645 2720 3649
rect 3115 3649 3119 3653
rect 3123 3649 3127 3653
rect 3139 3645 3143 3649
rect 3154 3645 3158 3649
rect 3196 3649 3200 3653
rect 3204 3649 3208 3653
rect 3220 3645 3224 3649
rect 3235 3645 3239 3649
rect 3169 3641 3173 3645
rect 3177 3641 3181 3645
rect 2591 3636 2595 3640
rect 2599 3636 2603 3640
rect 2941 3636 2945 3640
rect 2949 3636 2953 3640
rect 2957 3636 2961 3640
rect 2965 3636 2969 3640
rect 2973 3636 2977 3640
rect 2981 3636 2985 3640
rect 2992 3636 2996 3640
rect 3009 3636 3013 3640
rect 3026 3636 3030 3640
rect 3035 3636 3039 3640
rect 3048 3636 3052 3640
rect 3056 3636 3060 3640
rect 3064 3636 3068 3640
rect 3081 3636 3085 3640
rect 3091 3636 3095 3640
rect 3099 3636 3103 3640
rect 3250 3641 3254 3645
rect 3258 3641 3262 3645
rect 1996 3590 2000 3594
rect 2004 3590 2008 3594
rect 2012 3590 2016 3594
rect 2020 3590 2024 3594
rect 2028 3590 2032 3594
rect 2036 3590 2040 3594
rect 2047 3590 2051 3594
rect 2064 3590 2068 3594
rect 2081 3590 2085 3594
rect 2090 3590 2094 3594
rect 2103 3590 2107 3594
rect 2111 3590 2115 3594
rect 2119 3590 2123 3594
rect 2136 3590 2140 3594
rect 2146 3590 2150 3594
rect 2154 3590 2158 3594
rect 1630 3580 1634 3584
rect 1638 3580 1642 3584
rect 1646 3580 1650 3584
rect 1659 3580 1663 3584
rect 1667 3580 1671 3584
rect 1675 3580 1679 3584
rect 1683 3580 1687 3584
rect 1691 3580 1695 3584
rect 1704 3580 1708 3584
rect 1717 3580 1721 3584
rect 1725 3580 1729 3584
rect 1733 3580 1737 3584
rect 1741 3580 1745 3584
rect 1754 3580 1758 3584
rect 2194 3589 2198 3593
rect 2209 3589 2213 3593
rect 2275 3589 2279 3593
rect 2290 3589 2294 3593
rect 2941 3590 2945 3594
rect 2949 3590 2953 3594
rect 2957 3590 2961 3594
rect 2965 3590 2969 3594
rect 2973 3590 2977 3594
rect 2981 3590 2985 3594
rect 2992 3590 2996 3594
rect 3009 3590 3013 3594
rect 3026 3590 3030 3594
rect 3035 3590 3039 3594
rect 3048 3590 3052 3594
rect 3056 3590 3060 3594
rect 3064 3590 3068 3594
rect 3081 3590 3085 3594
rect 3091 3590 3095 3594
rect 3099 3590 3103 3594
rect 2575 3580 2579 3584
rect 2583 3580 2587 3584
rect 2591 3580 2595 3584
rect 2604 3580 2608 3584
rect 2612 3580 2616 3584
rect 2620 3580 2624 3584
rect 2628 3580 2632 3584
rect 2636 3580 2640 3584
rect 2649 3580 2653 3584
rect 2662 3580 2666 3584
rect 2670 3580 2674 3584
rect 2678 3580 2682 3584
rect 2686 3580 2690 3584
rect 2699 3580 2703 3584
rect 3139 3589 3143 3593
rect 3154 3589 3158 3593
rect 3220 3589 3224 3593
rect 3235 3589 3239 3593
rect 2194 3513 2198 3517
rect 2209 3513 2213 3517
rect 2275 3517 2279 3521
rect 2283 3517 2287 3521
rect 2299 3513 2303 3517
rect 2314 3513 2318 3517
rect 2224 3509 2228 3513
rect 2232 3509 2236 3513
rect 1996 3504 2000 3508
rect 2004 3504 2008 3508
rect 2012 3504 2016 3508
rect 2020 3504 2024 3508
rect 2028 3504 2032 3508
rect 2036 3504 2040 3508
rect 2047 3504 2051 3508
rect 2064 3504 2068 3508
rect 2081 3504 2085 3508
rect 2090 3504 2094 3508
rect 2103 3504 2107 3508
rect 2111 3504 2115 3508
rect 2119 3504 2123 3508
rect 2136 3504 2140 3508
rect 2146 3504 2150 3508
rect 2154 3504 2158 3508
rect 2329 3509 2333 3513
rect 2337 3509 2341 3513
rect 3139 3513 3143 3517
rect 3154 3513 3158 3517
rect 3220 3517 3224 3521
rect 3228 3517 3232 3521
rect 3244 3513 3248 3517
rect 3259 3513 3263 3517
rect 3169 3509 3173 3513
rect 3177 3509 3181 3513
rect 2941 3504 2945 3508
rect 2949 3504 2953 3508
rect 2957 3504 2961 3508
rect 2965 3504 2969 3508
rect 2973 3504 2977 3508
rect 2981 3504 2985 3508
rect 2992 3504 2996 3508
rect 3009 3504 3013 3508
rect 3026 3504 3030 3508
rect 3035 3504 3039 3508
rect 3048 3504 3052 3508
rect 3056 3504 3060 3508
rect 3064 3504 3068 3508
rect 3081 3504 3085 3508
rect 3091 3504 3095 3508
rect 3099 3504 3103 3508
rect 3274 3509 3278 3513
rect 3282 3509 3286 3513
rect 1996 3458 2000 3462
rect 2004 3458 2008 3462
rect 2012 3458 2016 3462
rect 2020 3458 2024 3462
rect 2028 3458 2032 3462
rect 2036 3458 2040 3462
rect 2047 3458 2051 3462
rect 2064 3458 2068 3462
rect 2081 3458 2085 3462
rect 2090 3458 2094 3462
rect 2103 3458 2107 3462
rect 2111 3458 2115 3462
rect 2119 3458 2123 3462
rect 2136 3458 2140 3462
rect 2146 3458 2150 3462
rect 2154 3458 2158 3462
rect 2194 3458 2198 3462
rect 2209 3458 2213 3462
rect 2299 3458 2303 3462
rect 2314 3458 2318 3462
rect 2941 3458 2945 3462
rect 2949 3458 2953 3462
rect 2957 3458 2961 3462
rect 2965 3458 2969 3462
rect 2973 3458 2977 3462
rect 2981 3458 2985 3462
rect 2992 3458 2996 3462
rect 3009 3458 3013 3462
rect 3026 3458 3030 3462
rect 3035 3458 3039 3462
rect 3048 3458 3052 3462
rect 3056 3458 3060 3462
rect 3064 3458 3068 3462
rect 3081 3458 3085 3462
rect 3091 3458 3095 3462
rect 3099 3458 3103 3462
rect 3139 3458 3143 3462
rect 3154 3458 3158 3462
rect 3244 3458 3248 3462
rect 3259 3458 3263 3462
rect 2194 3381 2198 3385
rect 2209 3381 2213 3385
rect 2251 3385 2255 3389
rect 2259 3385 2263 3389
rect 2275 3381 2279 3385
rect 2290 3381 2294 3385
rect 2341 3385 2345 3389
rect 2349 3385 2353 3389
rect 2365 3381 2369 3385
rect 2380 3381 2384 3385
rect 2224 3377 2228 3381
rect 2232 3377 2236 3381
rect 1996 3372 2000 3376
rect 2004 3372 2008 3376
rect 2012 3372 2016 3376
rect 2020 3372 2024 3376
rect 2028 3372 2032 3376
rect 2036 3372 2040 3376
rect 2047 3372 2051 3376
rect 2064 3372 2068 3376
rect 2081 3372 2085 3376
rect 2090 3372 2094 3376
rect 2103 3372 2107 3376
rect 2111 3372 2115 3376
rect 2119 3372 2123 3376
rect 2136 3372 2140 3376
rect 2146 3372 2150 3376
rect 2154 3372 2158 3376
rect 2305 3377 2309 3381
rect 2313 3377 2317 3381
rect 2395 3377 2399 3381
rect 2403 3377 2407 3381
rect 3139 3381 3143 3385
rect 3154 3381 3158 3385
rect 3196 3385 3200 3389
rect 3204 3385 3208 3389
rect 3220 3381 3224 3385
rect 3235 3381 3239 3385
rect 3286 3385 3290 3389
rect 3294 3385 3298 3389
rect 3310 3381 3314 3385
rect 3325 3381 3329 3385
rect 3169 3377 3173 3381
rect 3177 3377 3181 3381
rect 2941 3372 2945 3376
rect 2949 3372 2953 3376
rect 2957 3372 2961 3376
rect 2965 3372 2969 3376
rect 2973 3372 2977 3376
rect 2981 3372 2985 3376
rect 2992 3372 2996 3376
rect 3009 3372 3013 3376
rect 3026 3372 3030 3376
rect 3035 3372 3039 3376
rect 3048 3372 3052 3376
rect 3056 3372 3060 3376
rect 3064 3372 3068 3376
rect 3081 3372 3085 3376
rect 3091 3372 3095 3376
rect 3099 3372 3103 3376
rect 3250 3377 3254 3381
rect 3258 3377 3262 3381
rect 3340 3377 3344 3381
rect 3348 3377 3352 3381
rect 1996 3326 2000 3330
rect 2004 3326 2008 3330
rect 2012 3326 2016 3330
rect 2020 3326 2024 3330
rect 2028 3326 2032 3330
rect 2036 3326 2040 3330
rect 2047 3326 2051 3330
rect 2064 3326 2068 3330
rect 2081 3326 2085 3330
rect 2090 3326 2094 3330
rect 2103 3326 2107 3330
rect 2111 3326 2115 3330
rect 2119 3326 2123 3330
rect 2136 3326 2140 3330
rect 2146 3326 2150 3330
rect 2154 3326 2158 3330
rect 2194 3323 2198 3327
rect 2209 3323 2213 3327
rect 2275 3323 2279 3327
rect 2290 3323 2294 3327
rect 2365 3323 2369 3327
rect 2380 3323 2384 3327
rect 2941 3326 2945 3330
rect 2949 3326 2953 3330
rect 2957 3326 2961 3330
rect 2965 3326 2969 3330
rect 2973 3326 2977 3330
rect 2981 3326 2985 3330
rect 2992 3326 2996 3330
rect 3009 3326 3013 3330
rect 3026 3326 3030 3330
rect 3035 3326 3039 3330
rect 3048 3326 3052 3330
rect 3056 3326 3060 3330
rect 3064 3326 3068 3330
rect 3081 3326 3085 3330
rect 3091 3326 3095 3330
rect 3099 3326 3103 3330
rect 3139 3323 3143 3327
rect 3154 3323 3158 3327
rect 3220 3323 3224 3327
rect 3235 3323 3239 3327
rect 3310 3323 3314 3327
rect 3325 3323 3329 3327
rect 2194 3249 2198 3253
rect 2209 3249 2213 3253
rect 2224 3245 2228 3249
rect 2232 3245 2236 3249
rect 1996 3240 2000 3244
rect 2004 3240 2008 3244
rect 2012 3240 2016 3244
rect 2020 3240 2024 3244
rect 2028 3240 2032 3244
rect 2036 3240 2040 3244
rect 2047 3240 2051 3244
rect 2064 3240 2068 3244
rect 2081 3240 2085 3244
rect 2090 3240 2094 3244
rect 2103 3240 2107 3244
rect 2111 3240 2115 3244
rect 2119 3240 2123 3244
rect 2136 3240 2140 3244
rect 2146 3240 2150 3244
rect 2154 3240 2158 3244
rect 3139 3249 3143 3253
rect 3154 3249 3158 3253
rect 3169 3245 3173 3249
rect 3177 3245 3181 3249
rect 2941 3240 2945 3244
rect 2949 3240 2953 3244
rect 2957 3240 2961 3244
rect 2965 3240 2969 3244
rect 2973 3240 2977 3244
rect 2981 3240 2985 3244
rect 2992 3240 2996 3244
rect 3009 3240 3013 3244
rect 3026 3240 3030 3244
rect 3035 3240 3039 3244
rect 3048 3240 3052 3244
rect 3056 3240 3060 3244
rect 3064 3240 3068 3244
rect 3081 3240 3085 3244
rect 3091 3240 3095 3244
rect 3099 3240 3103 3244
rect 1996 3194 2000 3198
rect 2004 3194 2008 3198
rect 2012 3194 2016 3198
rect 2020 3194 2024 3198
rect 2028 3194 2032 3198
rect 2036 3194 2040 3198
rect 2047 3194 2051 3198
rect 2064 3194 2068 3198
rect 2081 3194 2085 3198
rect 2090 3194 2094 3198
rect 2103 3194 2107 3198
rect 2111 3194 2115 3198
rect 2119 3194 2123 3198
rect 2136 3194 2140 3198
rect 2146 3194 2150 3198
rect 2154 3194 2158 3198
rect 2230 3194 2234 3198
rect 2238 3194 2242 3198
rect 2248 3194 2252 3198
rect 2256 3194 2260 3198
rect 2265 3194 2269 3198
rect 2273 3194 2277 3198
rect 2281 3194 2285 3198
rect 2289 3194 2293 3198
rect 2297 3194 2301 3198
rect 2308 3194 2312 3198
rect 2325 3194 2329 3198
rect 2342 3194 2346 3198
rect 2351 3194 2355 3198
rect 2364 3194 2368 3198
rect 2372 3194 2376 3198
rect 2380 3194 2384 3198
rect 2397 3194 2401 3198
rect 2407 3194 2411 3198
rect 2415 3194 2419 3198
rect 1507 3180 1511 3184
rect 1520 3180 1524 3184
rect 1528 3180 1532 3184
rect 1536 3180 1540 3184
rect 1544 3180 1548 3184
rect 1557 3180 1561 3184
rect 1570 3180 1574 3184
rect 1578 3180 1582 3184
rect 1586 3180 1590 3184
rect 1594 3180 1598 3184
rect 1602 3180 1606 3184
rect 1615 3180 1619 3184
rect 1623 3180 1627 3184
rect 1631 3180 1635 3184
rect 1639 3180 1643 3184
rect 1652 3180 1656 3184
rect 1660 3180 1664 3184
rect 1668 3180 1672 3184
rect 1676 3180 1680 3184
rect 1689 3180 1693 3184
rect 1702 3180 1706 3184
rect 1710 3180 1714 3184
rect 1718 3180 1722 3184
rect 1726 3180 1730 3184
rect 1734 3180 1738 3184
rect 1747 3180 1751 3184
rect 1755 3180 1759 3184
rect 1763 3180 1767 3184
rect 1771 3180 1775 3184
rect 1784 3180 1788 3184
rect 1792 3180 1796 3184
rect 1800 3180 1804 3184
rect 1808 3180 1812 3184
rect 1821 3180 1825 3184
rect 1834 3180 1838 3184
rect 1842 3180 1846 3184
rect 1850 3180 1854 3184
rect 1858 3180 1862 3184
rect 1866 3180 1870 3184
rect 1879 3180 1883 3184
rect 1887 3180 1891 3184
rect 1895 3180 1899 3184
rect 2194 3187 2198 3191
rect 2209 3187 2213 3191
rect 2941 3194 2945 3198
rect 2949 3194 2953 3198
rect 2957 3194 2961 3198
rect 2965 3194 2969 3198
rect 2973 3194 2977 3198
rect 2981 3194 2985 3198
rect 2992 3194 2996 3198
rect 3009 3194 3013 3198
rect 3026 3194 3030 3198
rect 3035 3194 3039 3198
rect 3048 3194 3052 3198
rect 3056 3194 3060 3198
rect 3064 3194 3068 3198
rect 3081 3194 3085 3198
rect 3091 3194 3095 3198
rect 3099 3194 3103 3198
rect 3175 3194 3179 3198
rect 3183 3194 3187 3198
rect 3193 3194 3197 3198
rect 3201 3194 3205 3198
rect 3210 3194 3214 3198
rect 3218 3194 3222 3198
rect 3226 3194 3230 3198
rect 3234 3194 3238 3198
rect 3242 3194 3246 3198
rect 3253 3194 3257 3198
rect 3270 3194 3274 3198
rect 3287 3194 3291 3198
rect 3296 3194 3300 3198
rect 3309 3194 3313 3198
rect 3317 3194 3321 3198
rect 3325 3194 3329 3198
rect 3342 3194 3346 3198
rect 3352 3194 3356 3198
rect 3360 3194 3364 3198
rect 2452 3180 2456 3184
rect 2465 3180 2469 3184
rect 2473 3180 2477 3184
rect 2481 3180 2485 3184
rect 2489 3180 2493 3184
rect 2502 3180 2506 3184
rect 2515 3180 2519 3184
rect 2523 3180 2527 3184
rect 2531 3180 2535 3184
rect 2539 3180 2543 3184
rect 2547 3180 2551 3184
rect 2560 3180 2564 3184
rect 2568 3180 2572 3184
rect 2576 3180 2580 3184
rect 2584 3180 2588 3184
rect 2597 3180 2601 3184
rect 2605 3180 2609 3184
rect 2613 3180 2617 3184
rect 2621 3180 2625 3184
rect 2634 3180 2638 3184
rect 2647 3180 2651 3184
rect 2655 3180 2659 3184
rect 2663 3180 2667 3184
rect 2671 3180 2675 3184
rect 2679 3180 2683 3184
rect 2692 3180 2696 3184
rect 2700 3180 2704 3184
rect 2708 3180 2712 3184
rect 2716 3180 2720 3184
rect 2729 3180 2733 3184
rect 2737 3180 2741 3184
rect 2745 3180 2749 3184
rect 2753 3180 2757 3184
rect 2766 3180 2770 3184
rect 2779 3180 2783 3184
rect 2787 3180 2791 3184
rect 2795 3180 2799 3184
rect 2803 3180 2807 3184
rect 2811 3180 2815 3184
rect 2824 3180 2828 3184
rect 2832 3180 2836 3184
rect 2840 3180 2844 3184
rect 3139 3187 3143 3191
rect 3154 3187 3158 3191
rect 1622 3136 1626 3140
rect 1630 3136 1634 3140
rect 1646 3136 1650 3140
rect 1654 3136 1658 3140
rect 2424 3141 2428 3145
rect 2424 3132 2428 3137
rect 2567 3136 2571 3140
rect 2575 3136 2579 3140
rect 2591 3136 2595 3140
rect 2599 3136 2603 3140
rect 3369 3141 3373 3145
rect 3369 3132 3373 3137
rect 1642 3123 1646 3127
rect 1650 3123 1654 3127
rect 2587 3123 2591 3127
rect 2595 3123 2599 3127
rect 1638 3112 1642 3116
rect 2583 3112 2587 3116
rect 1638 3104 1642 3108
rect 1622 3100 1626 3104
rect 1630 3100 1634 3104
rect 1646 3100 1650 3104
rect 1654 3100 1658 3104
rect 2583 3104 2587 3108
rect 2567 3100 2571 3104
rect 2575 3100 2579 3104
rect 2591 3100 2595 3104
rect 2599 3100 2603 3104
rect 2290 3068 2294 3072
rect 2303 3068 2307 3072
rect 2311 3068 2315 3072
rect 2319 3068 2323 3072
rect 2327 3068 2331 3072
rect 2340 3068 2344 3072
rect 2353 3068 2357 3072
rect 2361 3068 2365 3072
rect 2369 3068 2373 3072
rect 2377 3068 2381 3072
rect 2385 3068 2389 3072
rect 2398 3068 2402 3072
rect 2406 3068 2410 3072
rect 2414 3068 2418 3072
rect 3235 3068 3239 3072
rect 3248 3068 3252 3072
rect 3256 3068 3260 3072
rect 3264 3068 3268 3072
rect 3272 3068 3276 3072
rect 3285 3068 3289 3072
rect 3298 3068 3302 3072
rect 3306 3068 3310 3072
rect 3314 3068 3318 3072
rect 3322 3068 3326 3072
rect 3330 3068 3334 3072
rect 3343 3068 3347 3072
rect 3351 3068 3355 3072
rect 3359 3068 3363 3072
rect 1507 3038 1511 3042
rect 1520 3038 1524 3042
rect 1528 3038 1532 3042
rect 1536 3038 1540 3042
rect 1544 3038 1548 3042
rect 1557 3038 1561 3042
rect 1570 3038 1574 3042
rect 1578 3038 1582 3042
rect 1586 3038 1590 3042
rect 1594 3038 1598 3042
rect 1602 3038 1606 3042
rect 1615 3038 1619 3042
rect 1623 3038 1627 3042
rect 1631 3038 1635 3042
rect 1639 3038 1643 3042
rect 1652 3038 1656 3042
rect 1660 3038 1664 3042
rect 1668 3038 1672 3042
rect 1676 3038 1680 3042
rect 1689 3038 1693 3042
rect 1702 3038 1706 3042
rect 1710 3038 1714 3042
rect 1718 3038 1722 3042
rect 1726 3038 1730 3042
rect 1734 3038 1738 3042
rect 1747 3038 1751 3042
rect 1755 3038 1759 3042
rect 1763 3038 1767 3042
rect 1771 3038 1775 3042
rect 1784 3038 1788 3042
rect 1792 3038 1796 3042
rect 1800 3038 1804 3042
rect 1808 3038 1812 3042
rect 1821 3038 1825 3042
rect 1834 3038 1838 3042
rect 1842 3038 1846 3042
rect 1850 3038 1854 3042
rect 1858 3038 1862 3042
rect 1866 3038 1870 3042
rect 1879 3038 1883 3042
rect 1887 3038 1891 3042
rect 1895 3038 1899 3042
rect 2452 3038 2456 3042
rect 2465 3038 2469 3042
rect 2473 3038 2477 3042
rect 2481 3038 2485 3042
rect 2489 3038 2493 3042
rect 2502 3038 2506 3042
rect 2515 3038 2519 3042
rect 2523 3038 2527 3042
rect 2531 3038 2535 3042
rect 2539 3038 2543 3042
rect 2547 3038 2551 3042
rect 2560 3038 2564 3042
rect 2568 3038 2572 3042
rect 2576 3038 2580 3042
rect 2584 3038 2588 3042
rect 2597 3038 2601 3042
rect 2605 3038 2609 3042
rect 2613 3038 2617 3042
rect 2621 3038 2625 3042
rect 2634 3038 2638 3042
rect 2647 3038 2651 3042
rect 2655 3038 2659 3042
rect 2663 3038 2667 3042
rect 2671 3038 2675 3042
rect 2679 3038 2683 3042
rect 2692 3038 2696 3042
rect 2700 3038 2704 3042
rect 2708 3038 2712 3042
rect 2716 3038 2720 3042
rect 2729 3038 2733 3042
rect 2737 3038 2741 3042
rect 2745 3038 2749 3042
rect 2753 3038 2757 3042
rect 2766 3038 2770 3042
rect 2779 3038 2783 3042
rect 2787 3038 2791 3042
rect 2795 3038 2799 3042
rect 2803 3038 2807 3042
rect 2811 3038 2815 3042
rect 2824 3038 2828 3042
rect 2832 3038 2836 3042
rect 2840 3038 2844 3042
rect 2436 2995 2440 2999
rect 2436 2987 2440 2991
rect 3381 2995 3385 2999
rect 3381 2987 3385 2991
rect 2290 2982 2294 2986
rect 2303 2982 2307 2986
rect 2311 2982 2315 2986
rect 2319 2982 2323 2986
rect 2327 2982 2331 2986
rect 2340 2982 2344 2986
rect 2353 2982 2357 2986
rect 2361 2982 2365 2986
rect 2369 2982 2373 2986
rect 2377 2982 2381 2986
rect 2385 2982 2389 2986
rect 2398 2982 2402 2986
rect 2406 2982 2410 2986
rect 2414 2982 2418 2986
rect 3235 2982 3239 2986
rect 3248 2982 3252 2986
rect 3256 2982 3260 2986
rect 3264 2982 3268 2986
rect 3272 2982 3276 2986
rect 3285 2982 3289 2986
rect 3298 2982 3302 2986
rect 3306 2982 3310 2986
rect 3314 2982 3318 2986
rect 3322 2982 3326 2986
rect 3330 2982 3334 2986
rect 3343 2982 3347 2986
rect 3351 2982 3355 2986
rect 3359 2982 3363 2986
rect 1507 2952 1511 2956
rect 1520 2952 1524 2956
rect 1528 2952 1532 2956
rect 1536 2952 1540 2956
rect 1544 2952 1548 2956
rect 1557 2952 1561 2956
rect 1570 2952 1574 2956
rect 1578 2952 1582 2956
rect 1586 2952 1590 2956
rect 1594 2952 1598 2956
rect 1602 2952 1606 2956
rect 1615 2952 1619 2956
rect 1623 2952 1627 2956
rect 1631 2952 1635 2956
rect 1639 2952 1643 2956
rect 1652 2952 1656 2956
rect 1660 2952 1664 2956
rect 1668 2952 1672 2956
rect 1676 2952 1680 2956
rect 1689 2952 1693 2956
rect 1702 2952 1706 2956
rect 1710 2952 1714 2956
rect 1718 2952 1722 2956
rect 1726 2952 1730 2956
rect 1734 2952 1738 2956
rect 1747 2952 1751 2956
rect 1755 2952 1759 2956
rect 1763 2952 1767 2956
rect 1771 2952 1775 2956
rect 1784 2952 1788 2956
rect 1792 2952 1796 2956
rect 1800 2952 1804 2956
rect 1808 2952 1812 2956
rect 1821 2952 1825 2956
rect 1834 2952 1838 2956
rect 1842 2952 1846 2956
rect 1850 2952 1854 2956
rect 1858 2952 1862 2956
rect 1866 2952 1870 2956
rect 1879 2952 1883 2956
rect 1887 2952 1891 2956
rect 1895 2952 1899 2956
rect 2452 2952 2456 2956
rect 2465 2952 2469 2956
rect 2473 2952 2477 2956
rect 2481 2952 2485 2956
rect 2489 2952 2493 2956
rect 2502 2952 2506 2956
rect 2515 2952 2519 2956
rect 2523 2952 2527 2956
rect 2531 2952 2535 2956
rect 2539 2952 2543 2956
rect 2547 2952 2551 2956
rect 2560 2952 2564 2956
rect 2568 2952 2572 2956
rect 2576 2952 2580 2956
rect 2584 2952 2588 2956
rect 2597 2952 2601 2956
rect 2605 2952 2609 2956
rect 2613 2952 2617 2956
rect 2621 2952 2625 2956
rect 2634 2952 2638 2956
rect 2647 2952 2651 2956
rect 2655 2952 2659 2956
rect 2663 2952 2667 2956
rect 2671 2952 2675 2956
rect 2679 2952 2683 2956
rect 2692 2952 2696 2956
rect 2700 2952 2704 2956
rect 2708 2952 2712 2956
rect 2716 2952 2720 2956
rect 2729 2952 2733 2956
rect 2737 2952 2741 2956
rect 2745 2952 2749 2956
rect 2753 2952 2757 2956
rect 2766 2952 2770 2956
rect 2779 2952 2783 2956
rect 2787 2952 2791 2956
rect 2795 2952 2799 2956
rect 2803 2952 2807 2956
rect 2811 2952 2815 2956
rect 2824 2952 2828 2956
rect 2832 2952 2836 2956
rect 2840 2952 2844 2956
rect 1739 2908 1743 2912
rect 1747 2908 1751 2912
rect 1763 2908 1767 2912
rect 1771 2908 1775 2912
rect 2684 2908 2688 2912
rect 2692 2908 2696 2912
rect 2708 2908 2712 2912
rect 2716 2908 2720 2912
rect 1759 2897 1763 2901
rect 1767 2897 1771 2901
rect 2704 2897 2708 2901
rect 2712 2897 2716 2901
rect 1755 2886 1759 2890
rect 2700 2886 2704 2890
rect 1755 2878 1759 2882
rect 2700 2878 2704 2882
rect 1739 2874 1743 2878
rect 1747 2874 1751 2878
rect 1763 2874 1767 2878
rect 1771 2874 1775 2878
rect 2684 2874 2688 2878
rect 2692 2874 2696 2878
rect 2708 2874 2712 2878
rect 2716 2874 2720 2878
rect 1507 2812 1511 2816
rect 1520 2812 1524 2816
rect 1528 2812 1532 2816
rect 1536 2812 1540 2816
rect 1544 2812 1548 2816
rect 1557 2812 1561 2816
rect 1570 2812 1574 2816
rect 1578 2812 1582 2816
rect 1586 2812 1590 2816
rect 1594 2812 1598 2816
rect 1602 2812 1606 2816
rect 1615 2812 1619 2816
rect 1623 2812 1627 2816
rect 1631 2812 1635 2816
rect 1639 2812 1643 2816
rect 1652 2812 1656 2816
rect 1660 2812 1664 2816
rect 1668 2812 1672 2816
rect 1676 2812 1680 2816
rect 1689 2812 1693 2816
rect 1702 2812 1706 2816
rect 1710 2812 1714 2816
rect 1718 2812 1722 2816
rect 1726 2812 1730 2816
rect 1734 2812 1738 2816
rect 1747 2812 1751 2816
rect 1755 2812 1759 2816
rect 1763 2812 1767 2816
rect 1771 2812 1775 2816
rect 1784 2812 1788 2816
rect 1792 2812 1796 2816
rect 1800 2812 1804 2816
rect 1808 2812 1812 2816
rect 1821 2812 1825 2816
rect 1834 2812 1838 2816
rect 1842 2812 1846 2816
rect 1850 2812 1854 2816
rect 1858 2812 1862 2816
rect 1866 2812 1870 2816
rect 1879 2812 1883 2816
rect 1887 2812 1891 2816
rect 1895 2812 1899 2816
rect 2452 2812 2456 2816
rect 2465 2812 2469 2816
rect 2473 2812 2477 2816
rect 2481 2812 2485 2816
rect 2489 2812 2493 2816
rect 2502 2812 2506 2816
rect 2515 2812 2519 2816
rect 2523 2812 2527 2816
rect 2531 2812 2535 2816
rect 2539 2812 2543 2816
rect 2547 2812 2551 2816
rect 2560 2812 2564 2816
rect 2568 2812 2572 2816
rect 2576 2812 2580 2816
rect 2584 2812 2588 2816
rect 2597 2812 2601 2816
rect 2605 2812 2609 2816
rect 2613 2812 2617 2816
rect 2621 2812 2625 2816
rect 2634 2812 2638 2816
rect 2647 2812 2651 2816
rect 2655 2812 2659 2816
rect 2663 2812 2667 2816
rect 2671 2812 2675 2816
rect 2679 2812 2683 2816
rect 2692 2812 2696 2816
rect 2700 2812 2704 2816
rect 2708 2812 2712 2816
rect 2716 2812 2720 2816
rect 2729 2812 2733 2816
rect 2737 2812 2741 2816
rect 2745 2812 2749 2816
rect 2753 2812 2757 2816
rect 2766 2812 2770 2816
rect 2779 2812 2783 2816
rect 2787 2812 2791 2816
rect 2795 2812 2799 2816
rect 2803 2812 2807 2816
rect 2811 2812 2815 2816
rect 2824 2812 2828 2816
rect 2832 2812 2836 2816
rect 2840 2812 2844 2816
rect 1991 2733 1995 2737
rect 2004 2733 2008 2737
rect 2012 2733 2016 2737
rect 2020 2733 2024 2737
rect 2028 2733 2032 2737
rect 2041 2733 2045 2737
rect 2054 2733 2058 2737
rect 2062 2733 2066 2737
rect 2070 2733 2074 2737
rect 2078 2733 2082 2737
rect 2086 2733 2090 2737
rect 2099 2733 2103 2737
rect 2107 2733 2111 2737
rect 2115 2733 2119 2737
rect 2123 2733 2127 2737
rect 2136 2733 2140 2737
rect 2144 2733 2148 2737
rect 2152 2733 2156 2737
rect 2160 2733 2164 2737
rect 2173 2733 2177 2737
rect 2186 2733 2190 2737
rect 2194 2733 2198 2737
rect 2202 2733 2206 2737
rect 2210 2733 2214 2737
rect 2218 2733 2222 2737
rect 2231 2733 2235 2737
rect 2239 2733 2243 2737
rect 2247 2733 2251 2737
rect 2255 2733 2259 2737
rect 2268 2733 2272 2737
rect 2276 2733 2280 2737
rect 2284 2733 2288 2737
rect 2292 2733 2296 2737
rect 2305 2733 2309 2737
rect 2318 2733 2322 2737
rect 2326 2733 2330 2737
rect 2334 2733 2338 2737
rect 2342 2733 2346 2737
rect 2350 2733 2354 2737
rect 2363 2733 2367 2737
rect 2371 2733 2375 2737
rect 2379 2733 2383 2737
rect 2387 2733 2391 2737
rect 2400 2733 2404 2737
rect 2408 2733 2412 2737
rect 2416 2733 2420 2737
rect 2424 2733 2428 2737
rect 2437 2733 2441 2737
rect 2450 2733 2454 2737
rect 2458 2733 2462 2737
rect 2466 2733 2470 2737
rect 2474 2733 2478 2737
rect 2482 2733 2486 2737
rect 2495 2733 2499 2737
rect 2503 2733 2507 2737
rect 2511 2733 2515 2737
rect 2936 2733 2940 2737
rect 2949 2733 2953 2737
rect 2957 2733 2961 2737
rect 2965 2733 2969 2737
rect 2973 2733 2977 2737
rect 2986 2733 2990 2737
rect 2999 2733 3003 2737
rect 3007 2733 3011 2737
rect 3015 2733 3019 2737
rect 3023 2733 3027 2737
rect 3031 2733 3035 2737
rect 3044 2733 3048 2737
rect 3052 2733 3056 2737
rect 3060 2733 3064 2737
rect 3068 2733 3072 2737
rect 3081 2733 3085 2737
rect 3089 2733 3093 2737
rect 3097 2733 3101 2737
rect 3105 2733 3109 2737
rect 3118 2733 3122 2737
rect 3131 2733 3135 2737
rect 3139 2733 3143 2737
rect 3147 2733 3151 2737
rect 3155 2733 3159 2737
rect 3163 2733 3167 2737
rect 3176 2733 3180 2737
rect 3184 2733 3188 2737
rect 3192 2733 3196 2737
rect 3200 2733 3204 2737
rect 3213 2733 3217 2737
rect 3221 2733 3225 2737
rect 3229 2733 3233 2737
rect 3237 2733 3241 2737
rect 3250 2733 3254 2737
rect 3263 2733 3267 2737
rect 3271 2733 3275 2737
rect 3279 2733 3283 2737
rect 3287 2733 3291 2737
rect 3295 2733 3299 2737
rect 3308 2733 3312 2737
rect 3316 2733 3320 2737
rect 3324 2733 3328 2737
rect 3332 2733 3336 2737
rect 3345 2733 3349 2737
rect 3353 2733 3357 2737
rect 3361 2733 3365 2737
rect 3369 2733 3373 2737
rect 3382 2733 3386 2737
rect 3395 2733 3399 2737
rect 3403 2733 3407 2737
rect 3411 2733 3415 2737
rect 3419 2733 3423 2737
rect 3427 2733 3431 2737
rect 3440 2733 3444 2737
rect 3448 2733 3452 2737
rect 3456 2733 3460 2737
rect 1639 2700 1643 2704
rect 1652 2700 1656 2704
rect 1660 2700 1664 2704
rect 1668 2700 1672 2704
rect 1676 2700 1680 2704
rect 1689 2700 1693 2704
rect 1702 2700 1706 2704
rect 1710 2700 1714 2704
rect 1718 2700 1722 2704
rect 1726 2700 1730 2704
rect 1734 2700 1738 2704
rect 1747 2700 1751 2704
rect 1755 2700 1759 2704
rect 1763 2700 1767 2704
rect 2584 2700 2588 2704
rect 2597 2700 2601 2704
rect 2605 2700 2609 2704
rect 2613 2700 2617 2704
rect 2621 2700 2625 2704
rect 2634 2700 2638 2704
rect 2647 2700 2651 2704
rect 2655 2700 2659 2704
rect 2663 2700 2667 2704
rect 2671 2700 2675 2704
rect 2679 2700 2683 2704
rect 2692 2700 2696 2704
rect 2700 2700 2704 2704
rect 2708 2700 2712 2704
rect 1763 2663 1767 2667
rect 1771 2663 1775 2667
rect 2170 2667 2174 2671
rect 2178 2667 2182 2671
rect 2194 2663 2198 2667
rect 2209 2663 2213 2667
rect 2251 2667 2255 2671
rect 2259 2667 2263 2671
rect 2275 2663 2279 2667
rect 2290 2663 2294 2667
rect 2224 2659 2228 2663
rect 2232 2659 2236 2663
rect 1646 2654 1650 2658
rect 1654 2654 1658 2658
rect 1996 2654 2000 2658
rect 2004 2654 2008 2658
rect 2012 2654 2016 2658
rect 2020 2654 2024 2658
rect 2028 2654 2032 2658
rect 2036 2654 2040 2658
rect 2047 2654 2051 2658
rect 2064 2654 2068 2658
rect 2081 2654 2085 2658
rect 2090 2654 2094 2658
rect 2103 2654 2107 2658
rect 2111 2654 2115 2658
rect 2119 2654 2123 2658
rect 2136 2654 2140 2658
rect 2146 2654 2150 2658
rect 2154 2654 2158 2658
rect 2305 2659 2309 2663
rect 2313 2659 2317 2663
rect 2708 2663 2712 2667
rect 2716 2663 2720 2667
rect 3115 2667 3119 2671
rect 3123 2667 3127 2671
rect 3139 2663 3143 2667
rect 3154 2663 3158 2667
rect 3196 2667 3200 2671
rect 3204 2667 3208 2671
rect 3220 2663 3224 2667
rect 3235 2663 3239 2667
rect 3169 2659 3173 2663
rect 3177 2659 3181 2663
rect 2591 2654 2595 2658
rect 2599 2654 2603 2658
rect 2941 2654 2945 2658
rect 2949 2654 2953 2658
rect 2957 2654 2961 2658
rect 2965 2654 2969 2658
rect 2973 2654 2977 2658
rect 2981 2654 2985 2658
rect 2992 2654 2996 2658
rect 3009 2654 3013 2658
rect 3026 2654 3030 2658
rect 3035 2654 3039 2658
rect 3048 2654 3052 2658
rect 3056 2654 3060 2658
rect 3064 2654 3068 2658
rect 3081 2654 3085 2658
rect 3091 2654 3095 2658
rect 3099 2654 3103 2658
rect 3250 2659 3254 2663
rect 3258 2659 3262 2663
rect 1996 2608 2000 2612
rect 2004 2608 2008 2612
rect 2012 2608 2016 2612
rect 2020 2608 2024 2612
rect 2028 2608 2032 2612
rect 2036 2608 2040 2612
rect 2047 2608 2051 2612
rect 2064 2608 2068 2612
rect 2081 2608 2085 2612
rect 2090 2608 2094 2612
rect 2103 2608 2107 2612
rect 2111 2608 2115 2612
rect 2119 2608 2123 2612
rect 2136 2608 2140 2612
rect 2146 2608 2150 2612
rect 2154 2608 2158 2612
rect 1630 2598 1634 2602
rect 1638 2598 1642 2602
rect 1646 2598 1650 2602
rect 1659 2598 1663 2602
rect 1667 2598 1671 2602
rect 1675 2598 1679 2602
rect 1683 2598 1687 2602
rect 1691 2598 1695 2602
rect 1704 2598 1708 2602
rect 1717 2598 1721 2602
rect 1725 2598 1729 2602
rect 1733 2598 1737 2602
rect 1741 2598 1745 2602
rect 1754 2598 1758 2602
rect 2194 2607 2198 2611
rect 2209 2607 2213 2611
rect 2275 2607 2279 2611
rect 2290 2607 2294 2611
rect 2941 2608 2945 2612
rect 2949 2608 2953 2612
rect 2957 2608 2961 2612
rect 2965 2608 2969 2612
rect 2973 2608 2977 2612
rect 2981 2608 2985 2612
rect 2992 2608 2996 2612
rect 3009 2608 3013 2612
rect 3026 2608 3030 2612
rect 3035 2608 3039 2612
rect 3048 2608 3052 2612
rect 3056 2608 3060 2612
rect 3064 2608 3068 2612
rect 3081 2608 3085 2612
rect 3091 2608 3095 2612
rect 3099 2608 3103 2612
rect 2575 2598 2579 2602
rect 2583 2598 2587 2602
rect 2591 2598 2595 2602
rect 2604 2598 2608 2602
rect 2612 2598 2616 2602
rect 2620 2598 2624 2602
rect 2628 2598 2632 2602
rect 2636 2598 2640 2602
rect 2649 2598 2653 2602
rect 2662 2598 2666 2602
rect 2670 2598 2674 2602
rect 2678 2598 2682 2602
rect 2686 2598 2690 2602
rect 2699 2598 2703 2602
rect 3139 2607 3143 2611
rect 3154 2607 3158 2611
rect 3220 2607 3224 2611
rect 3235 2607 3239 2611
rect 2194 2531 2198 2535
rect 2209 2531 2213 2535
rect 2275 2535 2279 2539
rect 2283 2535 2287 2539
rect 2299 2531 2303 2535
rect 2314 2531 2318 2535
rect 2224 2527 2228 2531
rect 2232 2527 2236 2531
rect 1996 2522 2000 2526
rect 2004 2522 2008 2526
rect 2012 2522 2016 2526
rect 2020 2522 2024 2526
rect 2028 2522 2032 2526
rect 2036 2522 2040 2526
rect 2047 2522 2051 2526
rect 2064 2522 2068 2526
rect 2081 2522 2085 2526
rect 2090 2522 2094 2526
rect 2103 2522 2107 2526
rect 2111 2522 2115 2526
rect 2119 2522 2123 2526
rect 2136 2522 2140 2526
rect 2146 2522 2150 2526
rect 2154 2522 2158 2526
rect 2329 2527 2333 2531
rect 2337 2527 2341 2531
rect 3139 2531 3143 2535
rect 3154 2531 3158 2535
rect 3220 2535 3224 2539
rect 3228 2535 3232 2539
rect 3244 2531 3248 2535
rect 3259 2531 3263 2535
rect 3169 2527 3173 2531
rect 3177 2527 3181 2531
rect 2941 2522 2945 2526
rect 2949 2522 2953 2526
rect 2957 2522 2961 2526
rect 2965 2522 2969 2526
rect 2973 2522 2977 2526
rect 2981 2522 2985 2526
rect 2992 2522 2996 2526
rect 3009 2522 3013 2526
rect 3026 2522 3030 2526
rect 3035 2522 3039 2526
rect 3048 2522 3052 2526
rect 3056 2522 3060 2526
rect 3064 2522 3068 2526
rect 3081 2522 3085 2526
rect 3091 2522 3095 2526
rect 3099 2522 3103 2526
rect 3274 2527 3278 2531
rect 3282 2527 3286 2531
rect 1996 2476 2000 2480
rect 2004 2476 2008 2480
rect 2012 2476 2016 2480
rect 2020 2476 2024 2480
rect 2028 2476 2032 2480
rect 2036 2476 2040 2480
rect 2047 2476 2051 2480
rect 2064 2476 2068 2480
rect 2081 2476 2085 2480
rect 2090 2476 2094 2480
rect 2103 2476 2107 2480
rect 2111 2476 2115 2480
rect 2119 2476 2123 2480
rect 2136 2476 2140 2480
rect 2146 2476 2150 2480
rect 2154 2476 2158 2480
rect 2194 2476 2198 2480
rect 2209 2476 2213 2480
rect 2299 2476 2303 2480
rect 2314 2476 2318 2480
rect 2941 2476 2945 2480
rect 2949 2476 2953 2480
rect 2957 2476 2961 2480
rect 2965 2476 2969 2480
rect 2973 2476 2977 2480
rect 2981 2476 2985 2480
rect 2992 2476 2996 2480
rect 3009 2476 3013 2480
rect 3026 2476 3030 2480
rect 3035 2476 3039 2480
rect 3048 2476 3052 2480
rect 3056 2476 3060 2480
rect 3064 2476 3068 2480
rect 3081 2476 3085 2480
rect 3091 2476 3095 2480
rect 3099 2476 3103 2480
rect 3139 2476 3143 2480
rect 3154 2476 3158 2480
rect 3244 2476 3248 2480
rect 3259 2476 3263 2480
rect 2194 2399 2198 2403
rect 2209 2399 2213 2403
rect 2251 2403 2255 2407
rect 2259 2403 2263 2407
rect 2275 2399 2279 2403
rect 2290 2399 2294 2403
rect 2341 2403 2345 2407
rect 2349 2403 2353 2407
rect 2365 2399 2369 2403
rect 2380 2399 2384 2403
rect 2224 2395 2228 2399
rect 2232 2395 2236 2399
rect 1996 2390 2000 2394
rect 2004 2390 2008 2394
rect 2012 2390 2016 2394
rect 2020 2390 2024 2394
rect 2028 2390 2032 2394
rect 2036 2390 2040 2394
rect 2047 2390 2051 2394
rect 2064 2390 2068 2394
rect 2081 2390 2085 2394
rect 2090 2390 2094 2394
rect 2103 2390 2107 2394
rect 2111 2390 2115 2394
rect 2119 2390 2123 2394
rect 2136 2390 2140 2394
rect 2146 2390 2150 2394
rect 2154 2390 2158 2394
rect 2305 2395 2309 2399
rect 2313 2395 2317 2399
rect 2395 2395 2399 2399
rect 2403 2395 2407 2399
rect 3139 2399 3143 2403
rect 3154 2399 3158 2403
rect 3196 2403 3200 2407
rect 3204 2403 3208 2407
rect 3220 2399 3224 2403
rect 3235 2399 3239 2403
rect 3286 2403 3290 2407
rect 3294 2403 3298 2407
rect 3310 2399 3314 2403
rect 3325 2399 3329 2403
rect 3169 2395 3173 2399
rect 3177 2395 3181 2399
rect 2941 2390 2945 2394
rect 2949 2390 2953 2394
rect 2957 2390 2961 2394
rect 2965 2390 2969 2394
rect 2973 2390 2977 2394
rect 2981 2390 2985 2394
rect 2992 2390 2996 2394
rect 3009 2390 3013 2394
rect 3026 2390 3030 2394
rect 3035 2390 3039 2394
rect 3048 2390 3052 2394
rect 3056 2390 3060 2394
rect 3064 2390 3068 2394
rect 3081 2390 3085 2394
rect 3091 2390 3095 2394
rect 3099 2390 3103 2394
rect 3250 2395 3254 2399
rect 3258 2395 3262 2399
rect 3340 2395 3344 2399
rect 3348 2395 3352 2399
rect 1996 2344 2000 2348
rect 2004 2344 2008 2348
rect 2012 2344 2016 2348
rect 2020 2344 2024 2348
rect 2028 2344 2032 2348
rect 2036 2344 2040 2348
rect 2047 2344 2051 2348
rect 2064 2344 2068 2348
rect 2081 2344 2085 2348
rect 2090 2344 2094 2348
rect 2103 2344 2107 2348
rect 2111 2344 2115 2348
rect 2119 2344 2123 2348
rect 2136 2344 2140 2348
rect 2146 2344 2150 2348
rect 2154 2344 2158 2348
rect 2194 2341 2198 2345
rect 2209 2341 2213 2345
rect 2275 2341 2279 2345
rect 2290 2341 2294 2345
rect 2365 2341 2369 2345
rect 2380 2341 2384 2345
rect 2941 2344 2945 2348
rect 2949 2344 2953 2348
rect 2957 2344 2961 2348
rect 2965 2344 2969 2348
rect 2973 2344 2977 2348
rect 2981 2344 2985 2348
rect 2992 2344 2996 2348
rect 3009 2344 3013 2348
rect 3026 2344 3030 2348
rect 3035 2344 3039 2348
rect 3048 2344 3052 2348
rect 3056 2344 3060 2348
rect 3064 2344 3068 2348
rect 3081 2344 3085 2348
rect 3091 2344 3095 2348
rect 3099 2344 3103 2348
rect 3139 2341 3143 2345
rect 3154 2341 3158 2345
rect 3220 2341 3224 2345
rect 3235 2341 3239 2345
rect 3310 2341 3314 2345
rect 3325 2341 3329 2345
rect 2194 2267 2198 2271
rect 2209 2267 2213 2271
rect 2224 2263 2228 2267
rect 2232 2263 2236 2267
rect 1996 2258 2000 2262
rect 2004 2258 2008 2262
rect 2012 2258 2016 2262
rect 2020 2258 2024 2262
rect 2028 2258 2032 2262
rect 2036 2258 2040 2262
rect 2047 2258 2051 2262
rect 2064 2258 2068 2262
rect 2081 2258 2085 2262
rect 2090 2258 2094 2262
rect 2103 2258 2107 2262
rect 2111 2258 2115 2262
rect 2119 2258 2123 2262
rect 2136 2258 2140 2262
rect 2146 2258 2150 2262
rect 2154 2258 2158 2262
rect 3139 2267 3143 2271
rect 3154 2267 3158 2271
rect 3169 2263 3173 2267
rect 3177 2263 3181 2267
rect 2941 2258 2945 2262
rect 2949 2258 2953 2262
rect 2957 2258 2961 2262
rect 2965 2258 2969 2262
rect 2973 2258 2977 2262
rect 2981 2258 2985 2262
rect 2992 2258 2996 2262
rect 3009 2258 3013 2262
rect 3026 2258 3030 2262
rect 3035 2258 3039 2262
rect 3048 2258 3052 2262
rect 3056 2258 3060 2262
rect 3064 2258 3068 2262
rect 3081 2258 3085 2262
rect 3091 2258 3095 2262
rect 3099 2258 3103 2262
rect 1996 2212 2000 2216
rect 2004 2212 2008 2216
rect 2012 2212 2016 2216
rect 2020 2212 2024 2216
rect 2028 2212 2032 2216
rect 2036 2212 2040 2216
rect 2047 2212 2051 2216
rect 2064 2212 2068 2216
rect 2081 2212 2085 2216
rect 2090 2212 2094 2216
rect 2103 2212 2107 2216
rect 2111 2212 2115 2216
rect 2119 2212 2123 2216
rect 2136 2212 2140 2216
rect 2146 2212 2150 2216
rect 2154 2212 2158 2216
rect 2230 2212 2234 2216
rect 2238 2212 2242 2216
rect 2248 2212 2252 2216
rect 2256 2212 2260 2216
rect 2265 2212 2269 2216
rect 2273 2212 2277 2216
rect 2281 2212 2285 2216
rect 2289 2212 2293 2216
rect 2297 2212 2301 2216
rect 2308 2212 2312 2216
rect 2325 2212 2329 2216
rect 2342 2212 2346 2216
rect 2351 2212 2355 2216
rect 2364 2212 2368 2216
rect 2372 2212 2376 2216
rect 2380 2212 2384 2216
rect 2397 2212 2401 2216
rect 2407 2212 2411 2216
rect 2415 2212 2419 2216
rect 1507 2198 1511 2202
rect 1520 2198 1524 2202
rect 1528 2198 1532 2202
rect 1536 2198 1540 2202
rect 1544 2198 1548 2202
rect 1557 2198 1561 2202
rect 1570 2198 1574 2202
rect 1578 2198 1582 2202
rect 1586 2198 1590 2202
rect 1594 2198 1598 2202
rect 1602 2198 1606 2202
rect 1615 2198 1619 2202
rect 1623 2198 1627 2202
rect 1631 2198 1635 2202
rect 1639 2198 1643 2202
rect 1652 2198 1656 2202
rect 1660 2198 1664 2202
rect 1668 2198 1672 2202
rect 1676 2198 1680 2202
rect 1689 2198 1693 2202
rect 1702 2198 1706 2202
rect 1710 2198 1714 2202
rect 1718 2198 1722 2202
rect 1726 2198 1730 2202
rect 1734 2198 1738 2202
rect 1747 2198 1751 2202
rect 1755 2198 1759 2202
rect 1763 2198 1767 2202
rect 1771 2198 1775 2202
rect 1784 2198 1788 2202
rect 1792 2198 1796 2202
rect 1800 2198 1804 2202
rect 1808 2198 1812 2202
rect 1821 2198 1825 2202
rect 1834 2198 1838 2202
rect 1842 2198 1846 2202
rect 1850 2198 1854 2202
rect 1858 2198 1862 2202
rect 1866 2198 1870 2202
rect 1879 2198 1883 2202
rect 1887 2198 1891 2202
rect 1895 2198 1899 2202
rect 2194 2205 2198 2209
rect 2209 2205 2213 2209
rect 2941 2212 2945 2216
rect 2949 2212 2953 2216
rect 2957 2212 2961 2216
rect 2965 2212 2969 2216
rect 2973 2212 2977 2216
rect 2981 2212 2985 2216
rect 2992 2212 2996 2216
rect 3009 2212 3013 2216
rect 3026 2212 3030 2216
rect 3035 2212 3039 2216
rect 3048 2212 3052 2216
rect 3056 2212 3060 2216
rect 3064 2212 3068 2216
rect 3081 2212 3085 2216
rect 3091 2212 3095 2216
rect 3099 2212 3103 2216
rect 3175 2212 3179 2216
rect 3183 2212 3187 2216
rect 3193 2212 3197 2216
rect 3201 2212 3205 2216
rect 3210 2212 3214 2216
rect 3218 2212 3222 2216
rect 3226 2212 3230 2216
rect 3234 2212 3238 2216
rect 3242 2212 3246 2216
rect 3253 2212 3257 2216
rect 3270 2212 3274 2216
rect 3287 2212 3291 2216
rect 3296 2212 3300 2216
rect 3309 2212 3313 2216
rect 3317 2212 3321 2216
rect 3325 2212 3329 2216
rect 3342 2212 3346 2216
rect 3352 2212 3356 2216
rect 3360 2212 3364 2216
rect 2452 2198 2456 2202
rect 2465 2198 2469 2202
rect 2473 2198 2477 2202
rect 2481 2198 2485 2202
rect 2489 2198 2493 2202
rect 2502 2198 2506 2202
rect 2515 2198 2519 2202
rect 2523 2198 2527 2202
rect 2531 2198 2535 2202
rect 2539 2198 2543 2202
rect 2547 2198 2551 2202
rect 2560 2198 2564 2202
rect 2568 2198 2572 2202
rect 2576 2198 2580 2202
rect 2584 2198 2588 2202
rect 2597 2198 2601 2202
rect 2605 2198 2609 2202
rect 2613 2198 2617 2202
rect 2621 2198 2625 2202
rect 2634 2198 2638 2202
rect 2647 2198 2651 2202
rect 2655 2198 2659 2202
rect 2663 2198 2667 2202
rect 2671 2198 2675 2202
rect 2679 2198 2683 2202
rect 2692 2198 2696 2202
rect 2700 2198 2704 2202
rect 2708 2198 2712 2202
rect 2716 2198 2720 2202
rect 2729 2198 2733 2202
rect 2737 2198 2741 2202
rect 2745 2198 2749 2202
rect 2753 2198 2757 2202
rect 2766 2198 2770 2202
rect 2779 2198 2783 2202
rect 2787 2198 2791 2202
rect 2795 2198 2799 2202
rect 2803 2198 2807 2202
rect 2811 2198 2815 2202
rect 2824 2198 2828 2202
rect 2832 2198 2836 2202
rect 2840 2198 2844 2202
rect 3139 2205 3143 2209
rect 3154 2205 3158 2209
rect 1622 2154 1626 2158
rect 1630 2154 1634 2158
rect 1646 2154 1650 2158
rect 1654 2154 1658 2158
rect 2424 2159 2428 2163
rect 2424 2151 2428 2155
rect 2567 2154 2571 2158
rect 2575 2154 2579 2158
rect 2591 2154 2595 2158
rect 2599 2154 2603 2158
rect 3369 2159 3373 2163
rect 3369 2151 3373 2155
rect 1642 2141 1646 2145
rect 1650 2141 1654 2145
rect 2587 2141 2591 2145
rect 2595 2141 2599 2145
rect 1638 2130 1642 2134
rect 2583 2130 2587 2134
rect 1638 2122 1642 2126
rect 1622 2118 1626 2122
rect 1630 2118 1634 2122
rect 1646 2118 1650 2122
rect 1654 2118 1658 2122
rect 2583 2122 2587 2126
rect 2567 2118 2571 2122
rect 2575 2118 2579 2122
rect 2591 2118 2595 2122
rect 2599 2118 2603 2122
rect 2290 2086 2294 2090
rect 2303 2086 2307 2090
rect 2311 2086 2315 2090
rect 2319 2086 2323 2090
rect 2327 2086 2331 2090
rect 2340 2086 2344 2090
rect 2353 2086 2357 2090
rect 2361 2086 2365 2090
rect 2369 2086 2373 2090
rect 2377 2086 2381 2090
rect 2385 2086 2389 2090
rect 2398 2086 2402 2090
rect 2406 2086 2410 2090
rect 2414 2086 2418 2090
rect 3235 2086 3239 2090
rect 3248 2086 3252 2090
rect 3256 2086 3260 2090
rect 3264 2086 3268 2090
rect 3272 2086 3276 2090
rect 3285 2086 3289 2090
rect 3298 2086 3302 2090
rect 3306 2086 3310 2090
rect 3314 2086 3318 2090
rect 3322 2086 3326 2090
rect 3330 2086 3334 2090
rect 3343 2086 3347 2090
rect 3351 2086 3355 2090
rect 3359 2086 3363 2090
rect 1507 2056 1511 2060
rect 1520 2056 1524 2060
rect 1528 2056 1532 2060
rect 1536 2056 1540 2060
rect 1544 2056 1548 2060
rect 1557 2056 1561 2060
rect 1570 2056 1574 2060
rect 1578 2056 1582 2060
rect 1586 2056 1590 2060
rect 1594 2056 1598 2060
rect 1602 2056 1606 2060
rect 1615 2056 1619 2060
rect 1623 2056 1627 2060
rect 1631 2056 1635 2060
rect 1639 2056 1643 2060
rect 1652 2056 1656 2060
rect 1660 2056 1664 2060
rect 1668 2056 1672 2060
rect 1676 2056 1680 2060
rect 1689 2056 1693 2060
rect 1702 2056 1706 2060
rect 1710 2056 1714 2060
rect 1718 2056 1722 2060
rect 1726 2056 1730 2060
rect 1734 2056 1738 2060
rect 1747 2056 1751 2060
rect 1755 2056 1759 2060
rect 1763 2056 1767 2060
rect 1771 2056 1775 2060
rect 1784 2056 1788 2060
rect 1792 2056 1796 2060
rect 1800 2056 1804 2060
rect 1808 2056 1812 2060
rect 1821 2056 1825 2060
rect 1834 2056 1838 2060
rect 1842 2056 1846 2060
rect 1850 2056 1854 2060
rect 1858 2056 1862 2060
rect 1866 2056 1870 2060
rect 1879 2056 1883 2060
rect 1887 2056 1891 2060
rect 1895 2056 1899 2060
rect 2452 2056 2456 2060
rect 2465 2056 2469 2060
rect 2473 2056 2477 2060
rect 2481 2056 2485 2060
rect 2489 2056 2493 2060
rect 2502 2056 2506 2060
rect 2515 2056 2519 2060
rect 2523 2056 2527 2060
rect 2531 2056 2535 2060
rect 2539 2056 2543 2060
rect 2547 2056 2551 2060
rect 2560 2056 2564 2060
rect 2568 2056 2572 2060
rect 2576 2056 2580 2060
rect 2584 2056 2588 2060
rect 2597 2056 2601 2060
rect 2605 2056 2609 2060
rect 2613 2056 2617 2060
rect 2621 2056 2625 2060
rect 2634 2056 2638 2060
rect 2647 2056 2651 2060
rect 2655 2056 2659 2060
rect 2663 2056 2667 2060
rect 2671 2056 2675 2060
rect 2679 2056 2683 2060
rect 2692 2056 2696 2060
rect 2700 2056 2704 2060
rect 2708 2056 2712 2060
rect 2716 2056 2720 2060
rect 2729 2056 2733 2060
rect 2737 2056 2741 2060
rect 2745 2056 2749 2060
rect 2753 2056 2757 2060
rect 2766 2056 2770 2060
rect 2779 2056 2783 2060
rect 2787 2056 2791 2060
rect 2795 2056 2799 2060
rect 2803 2056 2807 2060
rect 2811 2056 2815 2060
rect 2824 2056 2828 2060
rect 2832 2056 2836 2060
rect 2840 2056 2844 2060
rect 2436 2013 2440 2017
rect 2436 2005 2440 2009
rect 3381 2013 3385 2017
rect 3381 2005 3385 2009
rect 2290 2000 2294 2004
rect 2303 2000 2307 2004
rect 2311 2000 2315 2004
rect 2319 2000 2323 2004
rect 2327 2000 2331 2004
rect 2340 2000 2344 2004
rect 2353 2000 2357 2004
rect 2361 2000 2365 2004
rect 2369 2000 2373 2004
rect 2377 2000 2381 2004
rect 2385 2000 2389 2004
rect 2398 2000 2402 2004
rect 2406 2000 2410 2004
rect 2414 2000 2418 2004
rect 3235 2000 3239 2004
rect 3248 2000 3252 2004
rect 3256 2000 3260 2004
rect 3264 2000 3268 2004
rect 3272 2000 3276 2004
rect 3285 2000 3289 2004
rect 3298 2000 3302 2004
rect 3306 2000 3310 2004
rect 3314 2000 3318 2004
rect 3322 2000 3326 2004
rect 3330 2000 3334 2004
rect 3343 2000 3347 2004
rect 3351 2000 3355 2004
rect 3359 2000 3363 2004
rect 1507 1970 1511 1974
rect 1520 1970 1524 1974
rect 1528 1970 1532 1974
rect 1536 1970 1540 1974
rect 1544 1970 1548 1974
rect 1557 1970 1561 1974
rect 1570 1970 1574 1974
rect 1578 1970 1582 1974
rect 1586 1970 1590 1974
rect 1594 1970 1598 1974
rect 1602 1970 1606 1974
rect 1615 1970 1619 1974
rect 1623 1970 1627 1974
rect 1631 1970 1635 1974
rect 1639 1970 1643 1974
rect 1652 1970 1656 1974
rect 1660 1970 1664 1974
rect 1668 1970 1672 1974
rect 1676 1970 1680 1974
rect 1689 1970 1693 1974
rect 1702 1970 1706 1974
rect 1710 1970 1714 1974
rect 1718 1970 1722 1974
rect 1726 1970 1730 1974
rect 1734 1970 1738 1974
rect 1747 1970 1751 1974
rect 1755 1970 1759 1974
rect 1763 1970 1767 1974
rect 1771 1970 1775 1974
rect 1784 1970 1788 1974
rect 1792 1970 1796 1974
rect 1800 1970 1804 1974
rect 1808 1970 1812 1974
rect 1821 1970 1825 1974
rect 1834 1970 1838 1974
rect 1842 1970 1846 1974
rect 1850 1970 1854 1974
rect 1858 1970 1862 1974
rect 1866 1970 1870 1974
rect 1879 1970 1883 1974
rect 1887 1970 1891 1974
rect 1895 1970 1899 1974
rect 2452 1970 2456 1974
rect 2465 1970 2469 1974
rect 2473 1970 2477 1974
rect 2481 1970 2485 1974
rect 2489 1970 2493 1974
rect 2502 1970 2506 1974
rect 2515 1970 2519 1974
rect 2523 1970 2527 1974
rect 2531 1970 2535 1974
rect 2539 1970 2543 1974
rect 2547 1970 2551 1974
rect 2560 1970 2564 1974
rect 2568 1970 2572 1974
rect 2576 1970 2580 1974
rect 2584 1970 2588 1974
rect 2597 1970 2601 1974
rect 2605 1970 2609 1974
rect 2613 1970 2617 1974
rect 2621 1970 2625 1974
rect 2634 1970 2638 1974
rect 2647 1970 2651 1974
rect 2655 1970 2659 1974
rect 2663 1970 2667 1974
rect 2671 1970 2675 1974
rect 2679 1970 2683 1974
rect 2692 1970 2696 1974
rect 2700 1970 2704 1974
rect 2708 1970 2712 1974
rect 2716 1970 2720 1974
rect 2729 1970 2733 1974
rect 2737 1970 2741 1974
rect 2745 1970 2749 1974
rect 2753 1970 2757 1974
rect 2766 1970 2770 1974
rect 2779 1970 2783 1974
rect 2787 1970 2791 1974
rect 2795 1970 2799 1974
rect 2803 1970 2807 1974
rect 2811 1970 2815 1974
rect 2824 1970 2828 1974
rect 2832 1970 2836 1974
rect 2840 1970 2844 1974
rect 1739 1926 1743 1930
rect 1747 1926 1751 1930
rect 1763 1926 1767 1930
rect 1771 1926 1775 1930
rect 2684 1926 2688 1930
rect 2692 1926 2696 1930
rect 2708 1926 2712 1930
rect 2716 1926 2720 1930
rect 1759 1915 1763 1919
rect 1767 1915 1771 1919
rect 2704 1915 2708 1919
rect 2712 1915 2716 1919
rect 1755 1904 1759 1908
rect 2700 1904 2704 1908
rect 1755 1896 1759 1900
rect 2700 1896 2704 1900
rect 1739 1892 1743 1896
rect 1747 1892 1751 1896
rect 1763 1892 1767 1896
rect 1771 1892 1775 1896
rect 2684 1892 2688 1896
rect 2692 1892 2696 1896
rect 2708 1892 2712 1896
rect 2716 1892 2720 1896
rect 1507 1830 1511 1834
rect 1520 1830 1524 1834
rect 1528 1830 1532 1834
rect 1536 1830 1540 1834
rect 1544 1830 1548 1834
rect 1557 1830 1561 1834
rect 1570 1830 1574 1834
rect 1578 1830 1582 1834
rect 1586 1830 1590 1834
rect 1594 1830 1598 1834
rect 1602 1830 1606 1834
rect 1615 1830 1619 1834
rect 1623 1830 1627 1834
rect 1631 1830 1635 1834
rect 1639 1830 1643 1834
rect 1652 1830 1656 1834
rect 1660 1830 1664 1834
rect 1668 1830 1672 1834
rect 1676 1830 1680 1834
rect 1689 1830 1693 1834
rect 1702 1830 1706 1834
rect 1710 1830 1714 1834
rect 1718 1830 1722 1834
rect 1726 1830 1730 1834
rect 1734 1830 1738 1834
rect 1747 1830 1751 1834
rect 1755 1830 1759 1834
rect 1763 1830 1767 1834
rect 1771 1830 1775 1834
rect 1784 1830 1788 1834
rect 1792 1830 1796 1834
rect 1800 1830 1804 1834
rect 1808 1830 1812 1834
rect 1821 1830 1825 1834
rect 1834 1830 1838 1834
rect 1842 1830 1846 1834
rect 1850 1830 1854 1834
rect 1858 1830 1862 1834
rect 1866 1830 1870 1834
rect 1879 1830 1883 1834
rect 1887 1830 1891 1834
rect 1895 1830 1899 1834
rect 2452 1830 2456 1834
rect 2465 1830 2469 1834
rect 2473 1830 2477 1834
rect 2481 1830 2485 1834
rect 2489 1830 2493 1834
rect 2502 1830 2506 1834
rect 2515 1830 2519 1834
rect 2523 1830 2527 1834
rect 2531 1830 2535 1834
rect 2539 1830 2543 1834
rect 2547 1830 2551 1834
rect 2560 1830 2564 1834
rect 2568 1830 2572 1834
rect 2576 1830 2580 1834
rect 2584 1830 2588 1834
rect 2597 1830 2601 1834
rect 2605 1830 2609 1834
rect 2613 1830 2617 1834
rect 2621 1830 2625 1834
rect 2634 1830 2638 1834
rect 2647 1830 2651 1834
rect 2655 1830 2659 1834
rect 2663 1830 2667 1834
rect 2671 1830 2675 1834
rect 2679 1830 2683 1834
rect 2692 1830 2696 1834
rect 2700 1830 2704 1834
rect 2708 1830 2712 1834
rect 2716 1830 2720 1834
rect 2729 1830 2733 1834
rect 2737 1830 2741 1834
rect 2745 1830 2749 1834
rect 2753 1830 2757 1834
rect 2766 1830 2770 1834
rect 2779 1830 2783 1834
rect 2787 1830 2791 1834
rect 2795 1830 2799 1834
rect 2803 1830 2807 1834
rect 2811 1830 2815 1834
rect 2824 1830 2828 1834
rect 2832 1830 2836 1834
rect 2840 1830 2844 1834
<< pdcontact >>
rect 2696 4268 2700 4276
rect 2704 4268 2708 4276
rect 2720 4262 2724 4270
rect 2735 4262 2739 4270
rect 2750 4268 2754 4276
rect 2758 4268 2762 4276
rect 2870 4243 2886 4273
rect 2890 4243 2906 4273
rect 2923 4243 2939 4273
rect 2943 4243 2959 4273
rect 2720 4166 2724 4174
rect 2735 4166 2739 4174
rect 2674 4138 2678 4146
rect 2682 4138 2686 4146
rect 2696 4138 2700 4146
rect 2704 4138 2708 4146
rect 2720 4132 2724 4140
rect 2735 4132 2739 4140
rect 2750 4138 2754 4146
rect 2758 4138 2762 4146
rect 2776 4113 2792 4143
rect 2796 4113 2812 4143
rect 2829 4113 2845 4143
rect 2849 4113 2865 4143
rect 2720 4036 2724 4044
rect 2735 4036 2739 4044
rect 1991 3738 1995 3746
rect 2004 3738 2008 3746
rect 2012 3738 2016 3746
rect 2020 3742 2024 3746
rect 2028 3738 2032 3746
rect 2041 3738 2045 3746
rect 2054 3738 2058 3746
rect 2062 3738 2066 3746
rect 2070 3738 2074 3746
rect 2078 3742 2082 3746
rect 2086 3738 2090 3746
rect 2099 3738 2103 3746
rect 2107 3738 2111 3746
rect 2115 3738 2119 3746
rect 2123 3738 2127 3746
rect 2136 3738 2140 3746
rect 2144 3738 2148 3746
rect 2152 3742 2156 3746
rect 2160 3738 2164 3746
rect 2173 3738 2177 3746
rect 2186 3738 2190 3746
rect 2194 3738 2198 3746
rect 2202 3738 2206 3746
rect 2210 3742 2214 3746
rect 2218 3738 2222 3746
rect 2231 3738 2235 3746
rect 2239 3738 2243 3746
rect 2247 3738 2251 3746
rect 2255 3738 2259 3746
rect 2268 3738 2272 3746
rect 2276 3738 2280 3746
rect 2284 3742 2288 3746
rect 2292 3738 2296 3746
rect 2305 3738 2309 3746
rect 2318 3738 2322 3746
rect 2326 3738 2330 3746
rect 2334 3738 2338 3746
rect 2342 3742 2346 3746
rect 2350 3738 2354 3746
rect 2363 3738 2367 3746
rect 2371 3738 2375 3746
rect 2379 3738 2383 3746
rect 2387 3738 2391 3746
rect 2400 3738 2404 3746
rect 2408 3738 2412 3746
rect 2416 3742 2420 3746
rect 2424 3738 2428 3746
rect 2437 3738 2441 3746
rect 2450 3738 2454 3746
rect 2458 3738 2462 3746
rect 2466 3738 2470 3746
rect 2474 3742 2478 3746
rect 2482 3738 2486 3746
rect 2495 3738 2499 3746
rect 2503 3738 2507 3746
rect 2511 3738 2515 3746
rect 2936 3738 2940 3746
rect 2949 3738 2953 3746
rect 2957 3738 2961 3746
rect 2965 3742 2969 3746
rect 2973 3738 2977 3746
rect 2986 3738 2990 3746
rect 2999 3738 3003 3746
rect 3007 3738 3011 3746
rect 3015 3738 3019 3746
rect 3023 3742 3027 3746
rect 3031 3738 3035 3746
rect 3044 3738 3048 3746
rect 3052 3738 3056 3746
rect 3060 3738 3064 3746
rect 3068 3738 3072 3746
rect 3081 3738 3085 3746
rect 3089 3738 3093 3746
rect 3097 3742 3101 3746
rect 3105 3738 3109 3746
rect 3118 3738 3122 3746
rect 3131 3738 3135 3746
rect 3139 3738 3143 3746
rect 3147 3738 3151 3746
rect 3155 3742 3159 3746
rect 3163 3738 3167 3746
rect 3176 3738 3180 3746
rect 3184 3738 3188 3746
rect 3192 3738 3196 3746
rect 3200 3738 3204 3746
rect 3213 3738 3217 3746
rect 3221 3738 3225 3746
rect 3229 3742 3233 3746
rect 3237 3738 3241 3746
rect 3250 3738 3254 3746
rect 3263 3738 3267 3746
rect 3271 3738 3275 3746
rect 3279 3738 3283 3746
rect 3287 3742 3291 3746
rect 3295 3738 3299 3746
rect 3308 3738 3312 3746
rect 3316 3738 3320 3746
rect 3324 3738 3328 3746
rect 3332 3738 3336 3746
rect 3345 3738 3349 3746
rect 3353 3738 3357 3746
rect 3361 3742 3365 3746
rect 3369 3738 3373 3746
rect 3382 3738 3386 3746
rect 3395 3738 3399 3746
rect 3403 3738 3407 3746
rect 3411 3738 3415 3746
rect 3419 3742 3423 3746
rect 3427 3738 3431 3746
rect 3440 3738 3444 3746
rect 3448 3738 3452 3746
rect 3456 3738 3460 3746
rect 1639 3705 1643 3713
rect 1652 3705 1656 3713
rect 1660 3705 1664 3713
rect 1668 3709 1672 3713
rect 1676 3705 1680 3713
rect 1689 3705 1693 3713
rect 1702 3705 1706 3713
rect 1710 3705 1714 3713
rect 1718 3705 1722 3713
rect 1726 3709 1730 3713
rect 1734 3705 1738 3713
rect 1747 3705 1751 3713
rect 1755 3705 1759 3713
rect 1763 3705 1767 3713
rect 2584 3705 2588 3713
rect 2597 3705 2601 3713
rect 2605 3705 2609 3713
rect 2613 3709 2617 3713
rect 2621 3705 2625 3713
rect 2634 3705 2638 3713
rect 2647 3705 2651 3713
rect 2655 3705 2659 3713
rect 2663 3705 2667 3713
rect 2671 3709 2675 3713
rect 2679 3705 2683 3713
rect 2692 3705 2696 3713
rect 2700 3705 2704 3713
rect 2708 3705 2712 3713
rect 2170 3667 2174 3675
rect 2178 3667 2182 3675
rect 1996 3654 2000 3662
rect 2004 3654 2008 3662
rect 2012 3654 2016 3662
rect 2020 3654 2024 3662
rect 2028 3654 2032 3662
rect 2036 3654 2040 3662
rect 2047 3654 2051 3662
rect 2064 3654 2068 3662
rect 2081 3654 2085 3662
rect 2090 3654 2094 3662
rect 2103 3654 2107 3662
rect 2111 3654 2115 3662
rect 2119 3654 2123 3662
rect 2136 3654 2140 3662
rect 2146 3654 2150 3662
rect 2154 3654 2158 3662
rect 2194 3661 2198 3669
rect 2209 3661 2213 3669
rect 2224 3667 2228 3675
rect 2232 3667 2236 3675
rect 2251 3667 2255 3675
rect 2259 3667 2263 3675
rect 2275 3661 2279 3669
rect 2290 3661 2294 3669
rect 2305 3667 2309 3675
rect 2313 3667 2317 3675
rect 3115 3667 3119 3675
rect 3123 3667 3127 3675
rect 2941 3654 2945 3662
rect 2949 3654 2953 3662
rect 2957 3654 2961 3662
rect 2965 3654 2969 3662
rect 2973 3654 2977 3662
rect 2981 3654 2985 3662
rect 2992 3654 2996 3662
rect 3009 3654 3013 3662
rect 3026 3654 3030 3662
rect 3035 3654 3039 3662
rect 3048 3654 3052 3662
rect 3056 3654 3060 3662
rect 3064 3654 3068 3662
rect 3081 3654 3085 3662
rect 3091 3654 3095 3662
rect 3099 3654 3103 3662
rect 3139 3661 3143 3669
rect 3154 3661 3158 3669
rect 3169 3667 3173 3675
rect 3177 3667 3181 3675
rect 3196 3667 3200 3675
rect 3204 3667 3208 3675
rect 3220 3661 3224 3669
rect 3235 3661 3239 3669
rect 3250 3667 3254 3675
rect 3258 3667 3262 3675
rect 1630 3603 1634 3611
rect 1638 3603 1642 3611
rect 1646 3603 1650 3611
rect 1659 3603 1663 3611
rect 1667 3607 1671 3611
rect 1675 3603 1679 3611
rect 1683 3603 1687 3611
rect 1691 3603 1695 3611
rect 1704 3603 1708 3611
rect 1717 3603 1721 3611
rect 1725 3607 1729 3611
rect 1733 3603 1737 3611
rect 1741 3603 1745 3611
rect 1754 3603 1758 3611
rect 2575 3603 2579 3611
rect 2583 3603 2587 3611
rect 2591 3603 2595 3611
rect 2604 3603 2608 3611
rect 2612 3607 2616 3611
rect 2620 3603 2624 3611
rect 2628 3603 2632 3611
rect 2636 3603 2640 3611
rect 2649 3603 2653 3611
rect 2662 3603 2666 3611
rect 2670 3607 2674 3611
rect 2678 3603 2682 3611
rect 2686 3603 2690 3611
rect 2699 3603 2703 3611
rect 1996 3568 2000 3576
rect 2004 3568 2008 3576
rect 2012 3568 2016 3576
rect 2020 3568 2024 3576
rect 2028 3568 2032 3576
rect 2036 3568 2040 3576
rect 2047 3568 2051 3576
rect 2064 3568 2068 3576
rect 2081 3568 2085 3576
rect 2090 3568 2094 3576
rect 2103 3568 2107 3576
rect 2111 3568 2115 3576
rect 2119 3568 2123 3576
rect 2136 3568 2140 3576
rect 2146 3568 2150 3576
rect 2154 3568 2158 3576
rect 2194 3569 2198 3577
rect 2209 3569 2213 3577
rect 2275 3569 2279 3577
rect 2290 3569 2294 3577
rect 2941 3568 2945 3576
rect 2949 3568 2953 3576
rect 2957 3568 2961 3576
rect 2965 3568 2969 3576
rect 2973 3568 2977 3576
rect 2981 3568 2985 3576
rect 2992 3568 2996 3576
rect 3009 3568 3013 3576
rect 3026 3568 3030 3576
rect 3035 3568 3039 3576
rect 3048 3568 3052 3576
rect 3056 3568 3060 3576
rect 3064 3568 3068 3576
rect 3081 3568 3085 3576
rect 3091 3568 3095 3576
rect 3099 3568 3103 3576
rect 3139 3569 3143 3577
rect 3154 3569 3158 3577
rect 3220 3569 3224 3577
rect 3235 3569 3239 3577
rect 1996 3522 2000 3530
rect 2004 3522 2008 3530
rect 2012 3522 2016 3530
rect 2020 3522 2024 3530
rect 2028 3522 2032 3530
rect 2036 3522 2040 3530
rect 2047 3522 2051 3530
rect 2064 3522 2068 3530
rect 2081 3522 2085 3530
rect 2090 3522 2094 3530
rect 2103 3522 2107 3530
rect 2111 3522 2115 3530
rect 2119 3522 2123 3530
rect 2136 3522 2140 3530
rect 2146 3522 2150 3530
rect 2154 3522 2158 3530
rect 2194 3529 2198 3537
rect 2209 3529 2213 3537
rect 2224 3535 2228 3543
rect 2232 3535 2236 3543
rect 2275 3535 2279 3543
rect 2283 3535 2287 3543
rect 2299 3529 2303 3537
rect 2314 3529 2318 3537
rect 2329 3535 2333 3543
rect 2337 3535 2341 3543
rect 2941 3522 2945 3530
rect 2949 3522 2953 3530
rect 2957 3522 2961 3530
rect 2965 3522 2969 3530
rect 2973 3522 2977 3530
rect 2981 3522 2985 3530
rect 2992 3522 2996 3530
rect 3009 3522 3013 3530
rect 3026 3522 3030 3530
rect 3035 3522 3039 3530
rect 3048 3522 3052 3530
rect 3056 3522 3060 3530
rect 3064 3522 3068 3530
rect 3081 3522 3085 3530
rect 3091 3522 3095 3530
rect 3099 3522 3103 3530
rect 3139 3529 3143 3537
rect 3154 3529 3158 3537
rect 3169 3535 3173 3543
rect 3177 3535 3181 3543
rect 3220 3535 3224 3543
rect 3228 3535 3232 3543
rect 3244 3529 3248 3537
rect 3259 3529 3263 3537
rect 3274 3535 3278 3543
rect 3282 3535 3286 3543
rect 1996 3436 2000 3444
rect 2004 3436 2008 3444
rect 2012 3436 2016 3444
rect 2020 3436 2024 3444
rect 2028 3436 2032 3444
rect 2036 3436 2040 3444
rect 2047 3436 2051 3444
rect 2064 3436 2068 3444
rect 2081 3436 2085 3444
rect 2090 3436 2094 3444
rect 2103 3436 2107 3444
rect 2111 3436 2115 3444
rect 2119 3436 2123 3444
rect 2136 3436 2140 3444
rect 2146 3436 2150 3444
rect 2154 3436 2158 3444
rect 2194 3438 2198 3446
rect 2209 3438 2213 3446
rect 2299 3438 2303 3446
rect 2314 3438 2318 3446
rect 2941 3436 2945 3444
rect 2949 3436 2953 3444
rect 2957 3436 2961 3444
rect 2965 3436 2969 3444
rect 2973 3436 2977 3444
rect 2981 3436 2985 3444
rect 2992 3436 2996 3444
rect 3009 3436 3013 3444
rect 3026 3436 3030 3444
rect 3035 3436 3039 3444
rect 3048 3436 3052 3444
rect 3056 3436 3060 3444
rect 3064 3436 3068 3444
rect 3081 3436 3085 3444
rect 3091 3436 3095 3444
rect 3099 3436 3103 3444
rect 3139 3438 3143 3446
rect 3154 3438 3158 3446
rect 3244 3438 3248 3446
rect 3259 3438 3263 3446
rect 1996 3390 2000 3398
rect 2004 3390 2008 3398
rect 2012 3390 2016 3398
rect 2020 3390 2024 3398
rect 2028 3390 2032 3398
rect 2036 3390 2040 3398
rect 2047 3390 2051 3398
rect 2064 3390 2068 3398
rect 2081 3390 2085 3398
rect 2090 3390 2094 3398
rect 2103 3390 2107 3398
rect 2111 3390 2115 3398
rect 2119 3390 2123 3398
rect 2136 3390 2140 3398
rect 2146 3390 2150 3398
rect 2154 3390 2158 3398
rect 2194 3397 2198 3405
rect 2209 3397 2213 3405
rect 2224 3403 2228 3411
rect 2232 3403 2236 3411
rect 2251 3403 2255 3411
rect 2259 3403 2263 3411
rect 2275 3397 2279 3405
rect 2290 3397 2294 3405
rect 2305 3403 2309 3411
rect 2313 3403 2317 3411
rect 2341 3403 2345 3411
rect 2349 3403 2353 3411
rect 2365 3397 2369 3405
rect 2380 3397 2384 3405
rect 2395 3403 2399 3411
rect 2403 3403 2407 3411
rect 2941 3390 2945 3398
rect 2949 3390 2953 3398
rect 2957 3390 2961 3398
rect 2965 3390 2969 3398
rect 2973 3390 2977 3398
rect 2981 3390 2985 3398
rect 2992 3390 2996 3398
rect 3009 3390 3013 3398
rect 3026 3390 3030 3398
rect 3035 3390 3039 3398
rect 3048 3390 3052 3398
rect 3056 3390 3060 3398
rect 3064 3390 3068 3398
rect 3081 3390 3085 3398
rect 3091 3390 3095 3398
rect 3099 3390 3103 3398
rect 3139 3397 3143 3405
rect 3154 3397 3158 3405
rect 3169 3403 3173 3411
rect 3177 3403 3181 3411
rect 3196 3403 3200 3411
rect 3204 3403 3208 3411
rect 3220 3397 3224 3405
rect 3235 3397 3239 3405
rect 3250 3403 3254 3411
rect 3258 3403 3262 3411
rect 3286 3403 3290 3411
rect 3294 3403 3298 3411
rect 3310 3397 3314 3405
rect 3325 3397 3329 3405
rect 3340 3403 3344 3411
rect 3348 3403 3352 3411
rect 1996 3304 2000 3312
rect 2004 3304 2008 3312
rect 2012 3304 2016 3312
rect 2020 3304 2024 3312
rect 2028 3304 2032 3312
rect 2036 3304 2040 3312
rect 2047 3304 2051 3312
rect 2064 3304 2068 3312
rect 2081 3304 2085 3312
rect 2090 3304 2094 3312
rect 2103 3304 2107 3312
rect 2111 3304 2115 3312
rect 2119 3304 2123 3312
rect 2136 3304 2140 3312
rect 2146 3304 2150 3312
rect 2154 3304 2158 3312
rect 2194 3303 2198 3311
rect 2209 3303 2213 3311
rect 2275 3303 2279 3311
rect 2290 3303 2294 3311
rect 2365 3303 2369 3311
rect 2380 3303 2384 3311
rect 2941 3304 2945 3312
rect 2949 3304 2953 3312
rect 2957 3304 2961 3312
rect 2965 3304 2969 3312
rect 2973 3304 2977 3312
rect 2981 3304 2985 3312
rect 2992 3304 2996 3312
rect 3009 3304 3013 3312
rect 3026 3304 3030 3312
rect 3035 3304 3039 3312
rect 3048 3304 3052 3312
rect 3056 3304 3060 3312
rect 3064 3304 3068 3312
rect 3081 3304 3085 3312
rect 3091 3304 3095 3312
rect 3099 3304 3103 3312
rect 3139 3303 3143 3311
rect 3154 3303 3158 3311
rect 3220 3303 3224 3311
rect 3235 3303 3239 3311
rect 3310 3303 3314 3311
rect 3325 3303 3329 3311
rect 1996 3258 2000 3266
rect 2004 3258 2008 3266
rect 2012 3258 2016 3266
rect 2020 3258 2024 3266
rect 2028 3258 2032 3266
rect 2036 3258 2040 3266
rect 2047 3258 2051 3266
rect 2064 3258 2068 3266
rect 2081 3258 2085 3266
rect 2090 3258 2094 3266
rect 2103 3258 2107 3266
rect 2111 3258 2115 3266
rect 2119 3258 2123 3266
rect 2136 3258 2140 3266
rect 2146 3258 2150 3266
rect 2154 3258 2158 3266
rect 2194 3265 2198 3273
rect 2209 3265 2213 3273
rect 2224 3271 2228 3279
rect 2232 3271 2236 3279
rect 2941 3258 2945 3266
rect 2949 3258 2953 3266
rect 2957 3258 2961 3266
rect 2965 3258 2969 3266
rect 2973 3258 2977 3266
rect 2981 3258 2985 3266
rect 2992 3258 2996 3266
rect 3009 3258 3013 3266
rect 3026 3258 3030 3266
rect 3035 3258 3039 3266
rect 3048 3258 3052 3266
rect 3056 3258 3060 3266
rect 3064 3258 3068 3266
rect 3081 3258 3085 3266
rect 3091 3258 3095 3266
rect 3099 3258 3103 3266
rect 3139 3265 3143 3273
rect 3154 3265 3158 3273
rect 3169 3271 3173 3279
rect 3177 3271 3181 3279
rect 1507 3203 1511 3211
rect 1520 3203 1524 3211
rect 1528 3203 1532 3211
rect 1536 3207 1540 3211
rect 1544 3203 1548 3211
rect 1557 3203 1561 3211
rect 1570 3203 1574 3211
rect 1578 3203 1582 3211
rect 1586 3203 1590 3211
rect 1594 3207 1598 3211
rect 1602 3203 1606 3211
rect 1615 3203 1619 3211
rect 1623 3203 1627 3211
rect 1631 3203 1635 3211
rect 1639 3203 1643 3211
rect 1652 3203 1656 3211
rect 1660 3203 1664 3211
rect 1668 3207 1672 3211
rect 1676 3203 1680 3211
rect 1689 3203 1693 3211
rect 1702 3203 1706 3211
rect 1710 3203 1714 3211
rect 1718 3203 1722 3211
rect 1726 3207 1730 3211
rect 1734 3203 1738 3211
rect 1747 3203 1751 3211
rect 1755 3203 1759 3211
rect 1763 3203 1767 3211
rect 1771 3203 1775 3211
rect 1784 3203 1788 3211
rect 1792 3203 1796 3211
rect 1800 3207 1804 3211
rect 1808 3203 1812 3211
rect 1821 3203 1825 3211
rect 1834 3203 1838 3211
rect 1842 3203 1846 3211
rect 1850 3203 1854 3211
rect 1858 3207 1862 3211
rect 1866 3203 1870 3211
rect 1879 3203 1883 3211
rect 1887 3203 1891 3211
rect 1895 3203 1899 3211
rect 2452 3203 2456 3211
rect 2465 3203 2469 3211
rect 2473 3203 2477 3211
rect 2481 3207 2485 3211
rect 2489 3203 2493 3211
rect 2502 3203 2506 3211
rect 2515 3203 2519 3211
rect 2523 3203 2527 3211
rect 2531 3203 2535 3211
rect 2539 3207 2543 3211
rect 2547 3203 2551 3211
rect 2560 3203 2564 3211
rect 2568 3203 2572 3211
rect 2576 3203 2580 3211
rect 2584 3203 2588 3211
rect 2597 3203 2601 3211
rect 2605 3203 2609 3211
rect 2613 3207 2617 3211
rect 2621 3203 2625 3211
rect 2634 3203 2638 3211
rect 2647 3203 2651 3211
rect 2655 3203 2659 3211
rect 2663 3203 2667 3211
rect 2671 3207 2675 3211
rect 2679 3203 2683 3211
rect 2692 3203 2696 3211
rect 2700 3203 2704 3211
rect 2708 3203 2712 3211
rect 2716 3203 2720 3211
rect 2729 3203 2733 3211
rect 2737 3203 2741 3211
rect 2745 3207 2749 3211
rect 2753 3203 2757 3211
rect 2766 3203 2770 3211
rect 2779 3203 2783 3211
rect 2787 3203 2791 3211
rect 2795 3203 2799 3211
rect 2803 3207 2807 3211
rect 2811 3203 2815 3211
rect 2824 3203 2828 3211
rect 2832 3203 2836 3211
rect 2840 3203 2844 3211
rect 1996 3172 2000 3180
rect 2004 3172 2008 3180
rect 2012 3172 2016 3180
rect 2020 3172 2024 3180
rect 2028 3172 2032 3180
rect 2036 3172 2040 3180
rect 2047 3172 2051 3180
rect 2064 3172 2068 3180
rect 2081 3172 2085 3180
rect 2090 3172 2094 3180
rect 2103 3172 2107 3180
rect 2111 3172 2115 3180
rect 2119 3172 2123 3180
rect 2136 3172 2140 3180
rect 2146 3172 2150 3180
rect 2154 3172 2158 3180
rect 2194 3167 2198 3175
rect 2209 3167 2213 3175
rect 2230 3172 2234 3180
rect 2238 3172 2242 3180
rect 2248 3172 2252 3180
rect 2256 3172 2260 3180
rect 2265 3172 2269 3180
rect 2273 3172 2277 3180
rect 2281 3172 2285 3180
rect 2289 3172 2293 3180
rect 2297 3172 2301 3180
rect 2308 3172 2312 3180
rect 2325 3172 2329 3180
rect 2342 3172 2346 3180
rect 2351 3172 2355 3180
rect 2364 3172 2368 3180
rect 2372 3172 2376 3180
rect 2380 3172 2384 3180
rect 2397 3172 2401 3180
rect 2407 3172 2411 3180
rect 2415 3172 2419 3180
rect 2941 3172 2945 3180
rect 2949 3172 2953 3180
rect 2957 3172 2961 3180
rect 2965 3172 2969 3180
rect 2973 3172 2977 3180
rect 2981 3172 2985 3180
rect 2992 3172 2996 3180
rect 3009 3172 3013 3180
rect 3026 3172 3030 3180
rect 3035 3172 3039 3180
rect 3048 3172 3052 3180
rect 3056 3172 3060 3180
rect 3064 3172 3068 3180
rect 3081 3172 3085 3180
rect 3091 3172 3095 3180
rect 3099 3172 3103 3180
rect 3139 3167 3143 3175
rect 3154 3167 3158 3175
rect 3175 3172 3179 3180
rect 3183 3172 3187 3180
rect 3193 3172 3197 3180
rect 3201 3172 3205 3180
rect 3210 3172 3214 3180
rect 3218 3172 3222 3180
rect 3226 3172 3230 3180
rect 3234 3172 3238 3180
rect 3242 3172 3246 3180
rect 3253 3172 3257 3180
rect 3270 3172 3274 3180
rect 3287 3172 3291 3180
rect 3296 3172 3300 3180
rect 3309 3172 3313 3180
rect 3317 3172 3321 3180
rect 3325 3172 3329 3180
rect 3342 3172 3346 3180
rect 3352 3172 3356 3180
rect 3360 3172 3364 3180
rect 2290 3091 2294 3099
rect 2303 3091 2307 3099
rect 2311 3091 2315 3099
rect 2319 3095 2323 3099
rect 2327 3091 2331 3099
rect 2340 3091 2344 3099
rect 2353 3091 2357 3099
rect 2361 3091 2365 3099
rect 2369 3091 2373 3099
rect 2377 3095 2381 3099
rect 2385 3091 2389 3099
rect 2398 3091 2402 3099
rect 2406 3091 2410 3099
rect 2414 3091 2418 3099
rect 3235 3091 3239 3099
rect 3248 3091 3252 3099
rect 3256 3091 3260 3099
rect 3264 3095 3268 3099
rect 3272 3091 3276 3099
rect 3285 3091 3289 3099
rect 3298 3091 3302 3099
rect 3306 3091 3310 3099
rect 3314 3091 3318 3099
rect 3322 3095 3326 3099
rect 3330 3091 3334 3099
rect 3343 3091 3347 3099
rect 3351 3091 3355 3099
rect 3359 3091 3363 3099
rect 1507 3061 1511 3069
rect 1520 3061 1524 3069
rect 1528 3061 1532 3069
rect 1536 3065 1540 3069
rect 1544 3061 1548 3069
rect 1557 3061 1561 3069
rect 1570 3061 1574 3069
rect 1578 3061 1582 3069
rect 1586 3061 1590 3069
rect 1594 3065 1598 3069
rect 1602 3061 1606 3069
rect 1615 3061 1619 3069
rect 1623 3061 1627 3069
rect 1631 3061 1635 3069
rect 1639 3061 1643 3069
rect 1652 3061 1656 3069
rect 1660 3061 1664 3069
rect 1668 3065 1672 3069
rect 1676 3061 1680 3069
rect 1689 3061 1693 3069
rect 1702 3061 1706 3069
rect 1710 3061 1714 3069
rect 1718 3061 1722 3069
rect 1726 3065 1730 3069
rect 1734 3061 1738 3069
rect 1747 3061 1751 3069
rect 1755 3061 1759 3069
rect 1763 3061 1767 3069
rect 1771 3061 1775 3069
rect 1784 3061 1788 3069
rect 1792 3061 1796 3069
rect 1800 3065 1804 3069
rect 1808 3061 1812 3069
rect 1821 3061 1825 3069
rect 1834 3061 1838 3069
rect 1842 3061 1846 3069
rect 1850 3061 1854 3069
rect 1858 3065 1862 3069
rect 1866 3061 1870 3069
rect 1879 3061 1883 3069
rect 1887 3061 1891 3069
rect 1895 3061 1899 3069
rect 2452 3061 2456 3069
rect 2465 3061 2469 3069
rect 2473 3061 2477 3069
rect 2481 3065 2485 3069
rect 2489 3061 2493 3069
rect 2502 3061 2506 3069
rect 2515 3061 2519 3069
rect 2523 3061 2527 3069
rect 2531 3061 2535 3069
rect 2539 3065 2543 3069
rect 2547 3061 2551 3069
rect 2560 3061 2564 3069
rect 2568 3061 2572 3069
rect 2576 3061 2580 3069
rect 2584 3061 2588 3069
rect 2597 3061 2601 3069
rect 2605 3061 2609 3069
rect 2613 3065 2617 3069
rect 2621 3061 2625 3069
rect 2634 3061 2638 3069
rect 2647 3061 2651 3069
rect 2655 3061 2659 3069
rect 2663 3061 2667 3069
rect 2671 3065 2675 3069
rect 2679 3061 2683 3069
rect 2692 3061 2696 3069
rect 2700 3061 2704 3069
rect 2708 3061 2712 3069
rect 2716 3061 2720 3069
rect 2729 3061 2733 3069
rect 2737 3061 2741 3069
rect 2745 3065 2749 3069
rect 2753 3061 2757 3069
rect 2766 3061 2770 3069
rect 2779 3061 2783 3069
rect 2787 3061 2791 3069
rect 2795 3061 2799 3069
rect 2803 3065 2807 3069
rect 2811 3061 2815 3069
rect 2824 3061 2828 3069
rect 2832 3061 2836 3069
rect 2840 3061 2844 3069
rect 2290 3005 2294 3013
rect 2303 3005 2307 3013
rect 2311 3005 2315 3013
rect 2319 3009 2323 3013
rect 2327 3005 2331 3013
rect 2340 3005 2344 3013
rect 2353 3005 2357 3013
rect 2361 3005 2365 3013
rect 2369 3005 2373 3013
rect 2377 3009 2381 3013
rect 2385 3005 2389 3013
rect 2398 3005 2402 3013
rect 2406 3005 2410 3013
rect 2414 3005 2418 3013
rect 3235 3005 3239 3013
rect 3248 3005 3252 3013
rect 3256 3005 3260 3013
rect 3264 3009 3268 3013
rect 3272 3005 3276 3013
rect 3285 3005 3289 3013
rect 3298 3005 3302 3013
rect 3306 3005 3310 3013
rect 3314 3005 3318 3013
rect 3322 3009 3326 3013
rect 3330 3005 3334 3013
rect 3343 3005 3347 3013
rect 3351 3005 3355 3013
rect 3359 3005 3363 3013
rect 1507 2975 1511 2983
rect 1520 2975 1524 2983
rect 1528 2975 1532 2983
rect 1536 2979 1540 2983
rect 1544 2975 1548 2983
rect 1557 2975 1561 2983
rect 1570 2975 1574 2983
rect 1578 2975 1582 2983
rect 1586 2975 1590 2983
rect 1594 2979 1598 2983
rect 1602 2975 1606 2983
rect 1615 2975 1619 2983
rect 1623 2975 1627 2983
rect 1631 2975 1635 2983
rect 1639 2975 1643 2983
rect 1652 2975 1656 2983
rect 1660 2975 1664 2983
rect 1668 2979 1672 2983
rect 1676 2975 1680 2983
rect 1689 2975 1693 2983
rect 1702 2975 1706 2983
rect 1710 2975 1714 2983
rect 1718 2975 1722 2983
rect 1726 2979 1730 2983
rect 1734 2975 1738 2983
rect 1747 2975 1751 2983
rect 1755 2975 1759 2983
rect 1763 2975 1767 2983
rect 1771 2975 1775 2983
rect 1784 2975 1788 2983
rect 1792 2975 1796 2983
rect 1800 2979 1804 2983
rect 1808 2975 1812 2983
rect 1821 2975 1825 2983
rect 1834 2975 1838 2983
rect 1842 2975 1846 2983
rect 1850 2975 1854 2983
rect 1858 2979 1862 2983
rect 1866 2975 1870 2983
rect 1879 2975 1883 2983
rect 1887 2975 1891 2983
rect 1895 2975 1899 2983
rect 2452 2975 2456 2983
rect 2465 2975 2469 2983
rect 2473 2975 2477 2983
rect 2481 2979 2485 2983
rect 2489 2975 2493 2983
rect 2502 2975 2506 2983
rect 2515 2975 2519 2983
rect 2523 2975 2527 2983
rect 2531 2975 2535 2983
rect 2539 2979 2543 2983
rect 2547 2975 2551 2983
rect 2560 2975 2564 2983
rect 2568 2975 2572 2983
rect 2576 2975 2580 2983
rect 2584 2975 2588 2983
rect 2597 2975 2601 2983
rect 2605 2975 2609 2983
rect 2613 2979 2617 2983
rect 2621 2975 2625 2983
rect 2634 2975 2638 2983
rect 2647 2975 2651 2983
rect 2655 2975 2659 2983
rect 2663 2975 2667 2983
rect 2671 2979 2675 2983
rect 2679 2975 2683 2983
rect 2692 2975 2696 2983
rect 2700 2975 2704 2983
rect 2708 2975 2712 2983
rect 2716 2975 2720 2983
rect 2729 2975 2733 2983
rect 2737 2975 2741 2983
rect 2745 2979 2749 2983
rect 2753 2975 2757 2983
rect 2766 2975 2770 2983
rect 2779 2975 2783 2983
rect 2787 2975 2791 2983
rect 2795 2975 2799 2983
rect 2803 2979 2807 2983
rect 2811 2975 2815 2983
rect 2824 2975 2828 2983
rect 2832 2975 2836 2983
rect 2840 2975 2844 2983
rect 1507 2835 1511 2843
rect 1520 2835 1524 2843
rect 1528 2835 1532 2843
rect 1536 2839 1540 2843
rect 1544 2835 1548 2843
rect 1557 2835 1561 2843
rect 1570 2835 1574 2843
rect 1578 2835 1582 2843
rect 1586 2835 1590 2843
rect 1594 2839 1598 2843
rect 1602 2835 1606 2843
rect 1615 2835 1619 2843
rect 1623 2835 1627 2843
rect 1631 2835 1635 2843
rect 1639 2835 1643 2843
rect 1652 2835 1656 2843
rect 1660 2835 1664 2843
rect 1668 2839 1672 2843
rect 1676 2835 1680 2843
rect 1689 2835 1693 2843
rect 1702 2835 1706 2843
rect 1710 2835 1714 2843
rect 1718 2835 1722 2843
rect 1726 2839 1730 2843
rect 1734 2835 1738 2843
rect 1747 2835 1751 2843
rect 1755 2835 1759 2843
rect 1763 2835 1767 2843
rect 1771 2835 1775 2843
rect 1784 2835 1788 2843
rect 1792 2835 1796 2843
rect 1800 2839 1804 2843
rect 1808 2835 1812 2843
rect 1821 2835 1825 2843
rect 1834 2835 1838 2843
rect 1842 2835 1846 2843
rect 1850 2835 1854 2843
rect 1858 2839 1862 2843
rect 1866 2835 1870 2843
rect 1879 2835 1883 2843
rect 1887 2835 1891 2843
rect 1895 2835 1899 2843
rect 2452 2835 2456 2843
rect 2465 2835 2469 2843
rect 2473 2835 2477 2843
rect 2481 2839 2485 2843
rect 2489 2835 2493 2843
rect 2502 2835 2506 2843
rect 2515 2835 2519 2843
rect 2523 2835 2527 2843
rect 2531 2835 2535 2843
rect 2539 2839 2543 2843
rect 2547 2835 2551 2843
rect 2560 2835 2564 2843
rect 2568 2835 2572 2843
rect 2576 2835 2580 2843
rect 2584 2835 2588 2843
rect 2597 2835 2601 2843
rect 2605 2835 2609 2843
rect 2613 2839 2617 2843
rect 2621 2835 2625 2843
rect 2634 2835 2638 2843
rect 2647 2835 2651 2843
rect 2655 2835 2659 2843
rect 2663 2835 2667 2843
rect 2671 2839 2675 2843
rect 2679 2835 2683 2843
rect 2692 2835 2696 2843
rect 2700 2835 2704 2843
rect 2708 2835 2712 2843
rect 2716 2835 2720 2843
rect 2729 2835 2733 2843
rect 2737 2835 2741 2843
rect 2745 2839 2749 2843
rect 2753 2835 2757 2843
rect 2766 2835 2770 2843
rect 2779 2835 2783 2843
rect 2787 2835 2791 2843
rect 2795 2835 2799 2843
rect 2803 2839 2807 2843
rect 2811 2835 2815 2843
rect 2824 2835 2828 2843
rect 2832 2835 2836 2843
rect 2840 2835 2844 2843
rect 1991 2756 1995 2764
rect 2004 2756 2008 2764
rect 2012 2756 2016 2764
rect 2020 2760 2024 2764
rect 2028 2756 2032 2764
rect 2041 2756 2045 2764
rect 2054 2756 2058 2764
rect 2062 2756 2066 2764
rect 2070 2756 2074 2764
rect 2078 2760 2082 2764
rect 2086 2756 2090 2764
rect 2099 2756 2103 2764
rect 2107 2756 2111 2764
rect 2115 2756 2119 2764
rect 2123 2756 2127 2764
rect 2136 2756 2140 2764
rect 2144 2756 2148 2764
rect 2152 2760 2156 2764
rect 2160 2756 2164 2764
rect 2173 2756 2177 2764
rect 2186 2756 2190 2764
rect 2194 2756 2198 2764
rect 2202 2756 2206 2764
rect 2210 2760 2214 2764
rect 2218 2756 2222 2764
rect 2231 2756 2235 2764
rect 2239 2756 2243 2764
rect 2247 2756 2251 2764
rect 2255 2756 2259 2764
rect 2268 2756 2272 2764
rect 2276 2756 2280 2764
rect 2284 2760 2288 2764
rect 2292 2756 2296 2764
rect 2305 2756 2309 2764
rect 2318 2756 2322 2764
rect 2326 2756 2330 2764
rect 2334 2756 2338 2764
rect 2342 2760 2346 2764
rect 2350 2756 2354 2764
rect 2363 2756 2367 2764
rect 2371 2756 2375 2764
rect 2379 2756 2383 2764
rect 2387 2756 2391 2764
rect 2400 2756 2404 2764
rect 2408 2756 2412 2764
rect 2416 2760 2420 2764
rect 2424 2756 2428 2764
rect 2437 2756 2441 2764
rect 2450 2756 2454 2764
rect 2458 2756 2462 2764
rect 2466 2756 2470 2764
rect 2474 2760 2478 2764
rect 2482 2756 2486 2764
rect 2495 2756 2499 2764
rect 2503 2756 2507 2764
rect 2511 2756 2515 2764
rect 2936 2756 2940 2764
rect 2949 2756 2953 2764
rect 2957 2756 2961 2764
rect 2965 2760 2969 2764
rect 2973 2756 2977 2764
rect 2986 2756 2990 2764
rect 2999 2756 3003 2764
rect 3007 2756 3011 2764
rect 3015 2756 3019 2764
rect 3023 2760 3027 2764
rect 3031 2756 3035 2764
rect 3044 2756 3048 2764
rect 3052 2756 3056 2764
rect 3060 2756 3064 2764
rect 3068 2756 3072 2764
rect 3081 2756 3085 2764
rect 3089 2756 3093 2764
rect 3097 2760 3101 2764
rect 3105 2756 3109 2764
rect 3118 2756 3122 2764
rect 3131 2756 3135 2764
rect 3139 2756 3143 2764
rect 3147 2756 3151 2764
rect 3155 2760 3159 2764
rect 3163 2756 3167 2764
rect 3176 2756 3180 2764
rect 3184 2756 3188 2764
rect 3192 2756 3196 2764
rect 3200 2756 3204 2764
rect 3213 2756 3217 2764
rect 3221 2756 3225 2764
rect 3229 2760 3233 2764
rect 3237 2756 3241 2764
rect 3250 2756 3254 2764
rect 3263 2756 3267 2764
rect 3271 2756 3275 2764
rect 3279 2756 3283 2764
rect 3287 2760 3291 2764
rect 3295 2756 3299 2764
rect 3308 2756 3312 2764
rect 3316 2756 3320 2764
rect 3324 2756 3328 2764
rect 3332 2756 3336 2764
rect 3345 2756 3349 2764
rect 3353 2756 3357 2764
rect 3361 2760 3365 2764
rect 3369 2756 3373 2764
rect 3382 2756 3386 2764
rect 3395 2756 3399 2764
rect 3403 2756 3407 2764
rect 3411 2756 3415 2764
rect 3419 2760 3423 2764
rect 3427 2756 3431 2764
rect 3440 2756 3444 2764
rect 3448 2756 3452 2764
rect 3456 2756 3460 2764
rect 1639 2723 1643 2731
rect 1652 2723 1656 2731
rect 1660 2723 1664 2731
rect 1668 2727 1672 2731
rect 1676 2723 1680 2731
rect 1689 2723 1693 2731
rect 1702 2723 1706 2731
rect 1710 2723 1714 2731
rect 1718 2723 1722 2731
rect 1726 2727 1730 2731
rect 1734 2723 1738 2731
rect 1747 2723 1751 2731
rect 1755 2723 1759 2731
rect 1763 2723 1767 2731
rect 2584 2723 2588 2731
rect 2597 2723 2601 2731
rect 2605 2723 2609 2731
rect 2613 2727 2617 2731
rect 2621 2723 2625 2731
rect 2634 2723 2638 2731
rect 2647 2723 2651 2731
rect 2655 2723 2659 2731
rect 2663 2723 2667 2731
rect 2671 2727 2675 2731
rect 2679 2723 2683 2731
rect 2692 2723 2696 2731
rect 2700 2723 2704 2731
rect 2708 2723 2712 2731
rect 2170 2685 2174 2693
rect 2178 2685 2182 2693
rect 1996 2672 2000 2680
rect 2004 2672 2008 2680
rect 2012 2672 2016 2680
rect 2020 2672 2024 2680
rect 2028 2672 2032 2680
rect 2036 2672 2040 2680
rect 2047 2672 2051 2680
rect 2064 2672 2068 2680
rect 2081 2672 2085 2680
rect 2090 2672 2094 2680
rect 2103 2672 2107 2680
rect 2111 2672 2115 2680
rect 2119 2672 2123 2680
rect 2136 2672 2140 2680
rect 2146 2672 2150 2680
rect 2154 2672 2158 2680
rect 2194 2679 2198 2687
rect 2209 2679 2213 2687
rect 2224 2685 2228 2693
rect 2232 2685 2236 2693
rect 2251 2685 2255 2693
rect 2259 2685 2263 2693
rect 2275 2679 2279 2687
rect 2290 2679 2294 2687
rect 2305 2685 2309 2693
rect 2313 2685 2317 2693
rect 3115 2685 3119 2693
rect 3123 2685 3127 2693
rect 2941 2672 2945 2680
rect 2949 2672 2953 2680
rect 2957 2672 2961 2680
rect 2965 2672 2969 2680
rect 2973 2672 2977 2680
rect 2981 2672 2985 2680
rect 2992 2672 2996 2680
rect 3009 2672 3013 2680
rect 3026 2672 3030 2680
rect 3035 2672 3039 2680
rect 3048 2672 3052 2680
rect 3056 2672 3060 2680
rect 3064 2672 3068 2680
rect 3081 2672 3085 2680
rect 3091 2672 3095 2680
rect 3099 2672 3103 2680
rect 3139 2679 3143 2687
rect 3154 2679 3158 2687
rect 3169 2685 3173 2693
rect 3177 2685 3181 2693
rect 3196 2685 3200 2693
rect 3204 2685 3208 2693
rect 3220 2679 3224 2687
rect 3235 2679 3239 2687
rect 3250 2685 3254 2693
rect 3258 2685 3262 2693
rect 1630 2621 1634 2629
rect 1638 2621 1642 2629
rect 1646 2621 1650 2629
rect 1659 2621 1663 2629
rect 1667 2625 1671 2629
rect 1675 2621 1679 2629
rect 1683 2621 1687 2629
rect 1691 2621 1695 2629
rect 1704 2621 1708 2629
rect 1717 2621 1721 2629
rect 1725 2625 1729 2629
rect 1733 2621 1737 2629
rect 1741 2621 1745 2629
rect 1754 2621 1758 2629
rect 2575 2621 2579 2629
rect 2583 2621 2587 2629
rect 2591 2621 2595 2629
rect 2604 2621 2608 2629
rect 2612 2625 2616 2629
rect 2620 2621 2624 2629
rect 2628 2621 2632 2629
rect 2636 2621 2640 2629
rect 2649 2621 2653 2629
rect 2662 2621 2666 2629
rect 2670 2625 2674 2629
rect 2678 2621 2682 2629
rect 2686 2621 2690 2629
rect 2699 2621 2703 2629
rect 1996 2586 2000 2594
rect 2004 2586 2008 2594
rect 2012 2586 2016 2594
rect 2020 2586 2024 2594
rect 2028 2586 2032 2594
rect 2036 2586 2040 2594
rect 2047 2586 2051 2594
rect 2064 2586 2068 2594
rect 2081 2586 2085 2594
rect 2090 2586 2094 2594
rect 2103 2586 2107 2594
rect 2111 2586 2115 2594
rect 2119 2586 2123 2594
rect 2136 2586 2140 2594
rect 2146 2586 2150 2594
rect 2154 2586 2158 2594
rect 2194 2587 2198 2595
rect 2209 2587 2213 2595
rect 2275 2587 2279 2595
rect 2290 2587 2294 2595
rect 2941 2586 2945 2594
rect 2949 2586 2953 2594
rect 2957 2586 2961 2594
rect 2965 2586 2969 2594
rect 2973 2586 2977 2594
rect 2981 2586 2985 2594
rect 2992 2586 2996 2594
rect 3009 2586 3013 2594
rect 3026 2586 3030 2594
rect 3035 2586 3039 2594
rect 3048 2586 3052 2594
rect 3056 2586 3060 2594
rect 3064 2586 3068 2594
rect 3081 2586 3085 2594
rect 3091 2586 3095 2594
rect 3099 2586 3103 2594
rect 3139 2587 3143 2595
rect 3154 2587 3158 2595
rect 3220 2587 3224 2595
rect 3235 2587 3239 2595
rect 1996 2540 2000 2548
rect 2004 2540 2008 2548
rect 2012 2540 2016 2548
rect 2020 2540 2024 2548
rect 2028 2540 2032 2548
rect 2036 2540 2040 2548
rect 2047 2540 2051 2548
rect 2064 2540 2068 2548
rect 2081 2540 2085 2548
rect 2090 2540 2094 2548
rect 2103 2540 2107 2548
rect 2111 2540 2115 2548
rect 2119 2540 2123 2548
rect 2136 2540 2140 2548
rect 2146 2540 2150 2548
rect 2154 2540 2158 2548
rect 2194 2547 2198 2555
rect 2209 2547 2213 2555
rect 2224 2553 2228 2561
rect 2232 2553 2236 2561
rect 2275 2553 2279 2561
rect 2283 2553 2287 2561
rect 2299 2547 2303 2555
rect 2314 2547 2318 2555
rect 2329 2553 2333 2561
rect 2337 2553 2341 2561
rect 2941 2540 2945 2548
rect 2949 2540 2953 2548
rect 2957 2540 2961 2548
rect 2965 2540 2969 2548
rect 2973 2540 2977 2548
rect 2981 2540 2985 2548
rect 2992 2540 2996 2548
rect 3009 2540 3013 2548
rect 3026 2540 3030 2548
rect 3035 2540 3039 2548
rect 3048 2540 3052 2548
rect 3056 2540 3060 2548
rect 3064 2540 3068 2548
rect 3081 2540 3085 2548
rect 3091 2540 3095 2548
rect 3099 2540 3103 2548
rect 3139 2547 3143 2555
rect 3154 2547 3158 2555
rect 3169 2553 3173 2561
rect 3177 2553 3181 2561
rect 3220 2553 3224 2561
rect 3228 2553 3232 2561
rect 3244 2547 3248 2555
rect 3259 2547 3263 2555
rect 3274 2553 3278 2561
rect 3282 2553 3286 2561
rect 1996 2454 2000 2462
rect 2004 2454 2008 2462
rect 2012 2454 2016 2462
rect 2020 2454 2024 2462
rect 2028 2454 2032 2462
rect 2036 2454 2040 2462
rect 2047 2454 2051 2462
rect 2064 2454 2068 2462
rect 2081 2454 2085 2462
rect 2090 2454 2094 2462
rect 2103 2454 2107 2462
rect 2111 2454 2115 2462
rect 2119 2454 2123 2462
rect 2136 2454 2140 2462
rect 2146 2454 2150 2462
rect 2154 2454 2158 2462
rect 2194 2456 2198 2464
rect 2209 2456 2213 2464
rect 2299 2456 2303 2464
rect 2314 2456 2318 2464
rect 2941 2454 2945 2462
rect 2949 2454 2953 2462
rect 2957 2454 2961 2462
rect 2965 2454 2969 2462
rect 2973 2454 2977 2462
rect 2981 2454 2985 2462
rect 2992 2454 2996 2462
rect 3009 2454 3013 2462
rect 3026 2454 3030 2462
rect 3035 2454 3039 2462
rect 3048 2454 3052 2462
rect 3056 2454 3060 2462
rect 3064 2454 3068 2462
rect 3081 2454 3085 2462
rect 3091 2454 3095 2462
rect 3099 2454 3103 2462
rect 3139 2456 3143 2464
rect 3154 2456 3158 2464
rect 3244 2456 3248 2464
rect 3259 2456 3263 2464
rect 1996 2408 2000 2416
rect 2004 2408 2008 2416
rect 2012 2408 2016 2416
rect 2020 2408 2024 2416
rect 2028 2408 2032 2416
rect 2036 2408 2040 2416
rect 2047 2408 2051 2416
rect 2064 2408 2068 2416
rect 2081 2408 2085 2416
rect 2090 2408 2094 2416
rect 2103 2408 2107 2416
rect 2111 2408 2115 2416
rect 2119 2408 2123 2416
rect 2136 2408 2140 2416
rect 2146 2408 2150 2416
rect 2154 2408 2158 2416
rect 2194 2415 2198 2423
rect 2209 2415 2213 2423
rect 2224 2421 2228 2429
rect 2232 2421 2236 2429
rect 2251 2421 2255 2429
rect 2259 2421 2263 2429
rect 2275 2415 2279 2423
rect 2290 2415 2294 2423
rect 2305 2421 2309 2429
rect 2313 2421 2317 2429
rect 2341 2421 2345 2429
rect 2349 2421 2353 2429
rect 2365 2415 2369 2423
rect 2380 2415 2384 2423
rect 2395 2421 2399 2429
rect 2403 2421 2407 2429
rect 2941 2408 2945 2416
rect 2949 2408 2953 2416
rect 2957 2408 2961 2416
rect 2965 2408 2969 2416
rect 2973 2408 2977 2416
rect 2981 2408 2985 2416
rect 2992 2408 2996 2416
rect 3009 2408 3013 2416
rect 3026 2408 3030 2416
rect 3035 2408 3039 2416
rect 3048 2408 3052 2416
rect 3056 2408 3060 2416
rect 3064 2408 3068 2416
rect 3081 2408 3085 2416
rect 3091 2408 3095 2416
rect 3099 2408 3103 2416
rect 3139 2415 3143 2423
rect 3154 2415 3158 2423
rect 3169 2421 3173 2429
rect 3177 2421 3181 2429
rect 3196 2421 3200 2429
rect 3204 2421 3208 2429
rect 3220 2415 3224 2423
rect 3235 2415 3239 2423
rect 3250 2421 3254 2429
rect 3258 2421 3262 2429
rect 3286 2421 3290 2429
rect 3294 2421 3298 2429
rect 3310 2415 3314 2423
rect 3325 2415 3329 2423
rect 3340 2421 3344 2429
rect 3348 2421 3352 2429
rect 1996 2322 2000 2330
rect 2004 2322 2008 2330
rect 2012 2322 2016 2330
rect 2020 2322 2024 2330
rect 2028 2322 2032 2330
rect 2036 2322 2040 2330
rect 2047 2322 2051 2330
rect 2064 2322 2068 2330
rect 2081 2322 2085 2330
rect 2090 2322 2094 2330
rect 2103 2322 2107 2330
rect 2111 2322 2115 2330
rect 2119 2322 2123 2330
rect 2136 2322 2140 2330
rect 2146 2322 2150 2330
rect 2154 2322 2158 2330
rect 2194 2321 2198 2329
rect 2209 2321 2213 2329
rect 2275 2321 2279 2329
rect 2290 2321 2294 2329
rect 2365 2321 2369 2329
rect 2380 2321 2384 2329
rect 2941 2322 2945 2330
rect 2949 2322 2953 2330
rect 2957 2322 2961 2330
rect 2965 2322 2969 2330
rect 2973 2322 2977 2330
rect 2981 2322 2985 2330
rect 2992 2322 2996 2330
rect 3009 2322 3013 2330
rect 3026 2322 3030 2330
rect 3035 2322 3039 2330
rect 3048 2322 3052 2330
rect 3056 2322 3060 2330
rect 3064 2322 3068 2330
rect 3081 2322 3085 2330
rect 3091 2322 3095 2330
rect 3099 2322 3103 2330
rect 3139 2321 3143 2329
rect 3154 2321 3158 2329
rect 3220 2321 3224 2329
rect 3235 2321 3239 2329
rect 3310 2321 3314 2329
rect 3325 2321 3329 2329
rect 1996 2276 2000 2284
rect 2004 2276 2008 2284
rect 2012 2276 2016 2284
rect 2020 2276 2024 2284
rect 2028 2276 2032 2284
rect 2036 2276 2040 2284
rect 2047 2276 2051 2284
rect 2064 2276 2068 2284
rect 2081 2276 2085 2284
rect 2090 2276 2094 2284
rect 2103 2276 2107 2284
rect 2111 2276 2115 2284
rect 2119 2276 2123 2284
rect 2136 2276 2140 2284
rect 2146 2276 2150 2284
rect 2154 2276 2158 2284
rect 2194 2283 2198 2291
rect 2209 2283 2213 2291
rect 2224 2289 2228 2297
rect 2232 2289 2236 2297
rect 2941 2276 2945 2284
rect 2949 2276 2953 2284
rect 2957 2276 2961 2284
rect 2965 2276 2969 2284
rect 2973 2276 2977 2284
rect 2981 2276 2985 2284
rect 2992 2276 2996 2284
rect 3009 2276 3013 2284
rect 3026 2276 3030 2284
rect 3035 2276 3039 2284
rect 3048 2276 3052 2284
rect 3056 2276 3060 2284
rect 3064 2276 3068 2284
rect 3081 2276 3085 2284
rect 3091 2276 3095 2284
rect 3099 2276 3103 2284
rect 3139 2283 3143 2291
rect 3154 2283 3158 2291
rect 3169 2289 3173 2297
rect 3177 2289 3181 2297
rect 1507 2221 1511 2229
rect 1520 2221 1524 2229
rect 1528 2221 1532 2229
rect 1536 2225 1540 2229
rect 1544 2221 1548 2229
rect 1557 2221 1561 2229
rect 1570 2221 1574 2229
rect 1578 2221 1582 2229
rect 1586 2221 1590 2229
rect 1594 2225 1598 2229
rect 1602 2221 1606 2229
rect 1615 2221 1619 2229
rect 1623 2221 1627 2229
rect 1631 2221 1635 2229
rect 1639 2221 1643 2229
rect 1652 2221 1656 2229
rect 1660 2221 1664 2229
rect 1668 2225 1672 2229
rect 1676 2221 1680 2229
rect 1689 2221 1693 2229
rect 1702 2221 1706 2229
rect 1710 2221 1714 2229
rect 1718 2221 1722 2229
rect 1726 2225 1730 2229
rect 1734 2221 1738 2229
rect 1747 2221 1751 2229
rect 1755 2221 1759 2229
rect 1763 2221 1767 2229
rect 1771 2221 1775 2229
rect 1784 2221 1788 2229
rect 1792 2221 1796 2229
rect 1800 2225 1804 2229
rect 1808 2221 1812 2229
rect 1821 2221 1825 2229
rect 1834 2221 1838 2229
rect 1842 2221 1846 2229
rect 1850 2221 1854 2229
rect 1858 2225 1862 2229
rect 1866 2221 1870 2229
rect 1879 2221 1883 2229
rect 1887 2221 1891 2229
rect 1895 2221 1899 2229
rect 2452 2221 2456 2229
rect 2465 2221 2469 2229
rect 2473 2221 2477 2229
rect 2481 2225 2485 2229
rect 2489 2221 2493 2229
rect 2502 2221 2506 2229
rect 2515 2221 2519 2229
rect 2523 2221 2527 2229
rect 2531 2221 2535 2229
rect 2539 2225 2543 2229
rect 2547 2221 2551 2229
rect 2560 2221 2564 2229
rect 2568 2221 2572 2229
rect 2576 2221 2580 2229
rect 2584 2221 2588 2229
rect 2597 2221 2601 2229
rect 2605 2221 2609 2229
rect 2613 2225 2617 2229
rect 2621 2221 2625 2229
rect 2634 2221 2638 2229
rect 2647 2221 2651 2229
rect 2655 2221 2659 2229
rect 2663 2221 2667 2229
rect 2671 2225 2675 2229
rect 2679 2221 2683 2229
rect 2692 2221 2696 2229
rect 2700 2221 2704 2229
rect 2708 2221 2712 2229
rect 2716 2221 2720 2229
rect 2729 2221 2733 2229
rect 2737 2221 2741 2229
rect 2745 2225 2749 2229
rect 2753 2221 2757 2229
rect 2766 2221 2770 2229
rect 2779 2221 2783 2229
rect 2787 2221 2791 2229
rect 2795 2221 2799 2229
rect 2803 2225 2807 2229
rect 2811 2221 2815 2229
rect 2824 2221 2828 2229
rect 2832 2221 2836 2229
rect 2840 2221 2844 2229
rect 1996 2190 2000 2198
rect 2004 2190 2008 2198
rect 2012 2190 2016 2198
rect 2020 2190 2024 2198
rect 2028 2190 2032 2198
rect 2036 2190 2040 2198
rect 2047 2190 2051 2198
rect 2064 2190 2068 2198
rect 2081 2190 2085 2198
rect 2090 2190 2094 2198
rect 2103 2190 2107 2198
rect 2111 2190 2115 2198
rect 2119 2190 2123 2198
rect 2136 2190 2140 2198
rect 2146 2190 2150 2198
rect 2154 2190 2158 2198
rect 2194 2185 2198 2193
rect 2209 2185 2213 2193
rect 2230 2190 2234 2198
rect 2238 2190 2242 2198
rect 2248 2190 2252 2198
rect 2256 2190 2260 2198
rect 2265 2190 2269 2198
rect 2273 2190 2277 2198
rect 2281 2190 2285 2198
rect 2289 2190 2293 2198
rect 2297 2190 2301 2198
rect 2308 2190 2312 2198
rect 2325 2190 2329 2198
rect 2342 2190 2346 2198
rect 2351 2190 2355 2198
rect 2364 2190 2368 2198
rect 2372 2190 2376 2198
rect 2380 2190 2384 2198
rect 2397 2190 2401 2198
rect 2407 2190 2411 2198
rect 2415 2190 2419 2198
rect 2941 2190 2945 2198
rect 2949 2190 2953 2198
rect 2957 2190 2961 2198
rect 2965 2190 2969 2198
rect 2973 2190 2977 2198
rect 2981 2190 2985 2198
rect 2992 2190 2996 2198
rect 3009 2190 3013 2198
rect 3026 2190 3030 2198
rect 3035 2190 3039 2198
rect 3048 2190 3052 2198
rect 3056 2190 3060 2198
rect 3064 2190 3068 2198
rect 3081 2190 3085 2198
rect 3091 2190 3095 2198
rect 3099 2190 3103 2198
rect 3139 2185 3143 2193
rect 3154 2185 3158 2193
rect 3175 2190 3179 2198
rect 3183 2190 3187 2198
rect 3193 2190 3197 2198
rect 3201 2190 3205 2198
rect 3210 2190 3214 2198
rect 3218 2190 3222 2198
rect 3226 2190 3230 2198
rect 3234 2190 3238 2198
rect 3242 2190 3246 2198
rect 3253 2190 3257 2198
rect 3270 2190 3274 2198
rect 3287 2190 3291 2198
rect 3296 2190 3300 2198
rect 3309 2190 3313 2198
rect 3317 2190 3321 2198
rect 3325 2190 3329 2198
rect 3342 2190 3346 2198
rect 3352 2190 3356 2198
rect 3360 2190 3364 2198
rect 2290 2109 2294 2117
rect 2303 2109 2307 2117
rect 2311 2109 2315 2117
rect 2319 2113 2323 2117
rect 2327 2109 2331 2117
rect 2340 2109 2344 2117
rect 2353 2109 2357 2117
rect 2361 2109 2365 2117
rect 2369 2109 2373 2117
rect 2377 2113 2381 2117
rect 2385 2109 2389 2117
rect 2398 2109 2402 2117
rect 2406 2109 2410 2117
rect 2414 2109 2418 2117
rect 3235 2109 3239 2117
rect 3248 2109 3252 2117
rect 3256 2109 3260 2117
rect 3264 2113 3268 2117
rect 3272 2109 3276 2117
rect 3285 2109 3289 2117
rect 3298 2109 3302 2117
rect 3306 2109 3310 2117
rect 3314 2109 3318 2117
rect 3322 2113 3326 2117
rect 3330 2109 3334 2117
rect 3343 2109 3347 2117
rect 3351 2109 3355 2117
rect 3359 2109 3363 2117
rect 1507 2079 1511 2087
rect 1520 2079 1524 2087
rect 1528 2079 1532 2087
rect 1536 2083 1540 2087
rect 1544 2079 1548 2087
rect 1557 2079 1561 2087
rect 1570 2079 1574 2087
rect 1578 2079 1582 2087
rect 1586 2079 1590 2087
rect 1594 2083 1598 2087
rect 1602 2079 1606 2087
rect 1615 2079 1619 2087
rect 1623 2079 1627 2087
rect 1631 2079 1635 2087
rect 1639 2079 1643 2087
rect 1652 2079 1656 2087
rect 1660 2079 1664 2087
rect 1668 2083 1672 2087
rect 1676 2079 1680 2087
rect 1689 2079 1693 2087
rect 1702 2079 1706 2087
rect 1710 2079 1714 2087
rect 1718 2079 1722 2087
rect 1726 2083 1730 2087
rect 1734 2079 1738 2087
rect 1747 2079 1751 2087
rect 1755 2079 1759 2087
rect 1763 2079 1767 2087
rect 1771 2079 1775 2087
rect 1784 2079 1788 2087
rect 1792 2079 1796 2087
rect 1800 2083 1804 2087
rect 1808 2079 1812 2087
rect 1821 2079 1825 2087
rect 1834 2079 1838 2087
rect 1842 2079 1846 2087
rect 1850 2079 1854 2087
rect 1858 2083 1862 2087
rect 1866 2079 1870 2087
rect 1879 2079 1883 2087
rect 1887 2079 1891 2087
rect 1895 2079 1899 2087
rect 2452 2079 2456 2087
rect 2465 2079 2469 2087
rect 2473 2079 2477 2087
rect 2481 2083 2485 2087
rect 2489 2079 2493 2087
rect 2502 2079 2506 2087
rect 2515 2079 2519 2087
rect 2523 2079 2527 2087
rect 2531 2079 2535 2087
rect 2539 2083 2543 2087
rect 2547 2079 2551 2087
rect 2560 2079 2564 2087
rect 2568 2079 2572 2087
rect 2576 2079 2580 2087
rect 2584 2079 2588 2087
rect 2597 2079 2601 2087
rect 2605 2079 2609 2087
rect 2613 2083 2617 2087
rect 2621 2079 2625 2087
rect 2634 2079 2638 2087
rect 2647 2079 2651 2087
rect 2655 2079 2659 2087
rect 2663 2079 2667 2087
rect 2671 2083 2675 2087
rect 2679 2079 2683 2087
rect 2692 2079 2696 2087
rect 2700 2079 2704 2087
rect 2708 2079 2712 2087
rect 2716 2079 2720 2087
rect 2729 2079 2733 2087
rect 2737 2079 2741 2087
rect 2745 2083 2749 2087
rect 2753 2079 2757 2087
rect 2766 2079 2770 2087
rect 2779 2079 2783 2087
rect 2787 2079 2791 2087
rect 2795 2079 2799 2087
rect 2803 2083 2807 2087
rect 2811 2079 2815 2087
rect 2824 2079 2828 2087
rect 2832 2079 2836 2087
rect 2840 2079 2844 2087
rect 2290 2023 2294 2031
rect 2303 2023 2307 2031
rect 2311 2023 2315 2031
rect 2319 2027 2323 2031
rect 2327 2023 2331 2031
rect 2340 2023 2344 2031
rect 2353 2023 2357 2031
rect 2361 2023 2365 2031
rect 2369 2023 2373 2031
rect 2377 2027 2381 2031
rect 2385 2023 2389 2031
rect 2398 2023 2402 2031
rect 2406 2023 2410 2031
rect 2414 2023 2418 2031
rect 3235 2023 3239 2031
rect 3248 2023 3252 2031
rect 3256 2023 3260 2031
rect 3264 2027 3268 2031
rect 3272 2023 3276 2031
rect 3285 2023 3289 2031
rect 3298 2023 3302 2031
rect 3306 2023 3310 2031
rect 3314 2023 3318 2031
rect 3322 2027 3326 2031
rect 3330 2023 3334 2031
rect 3343 2023 3347 2031
rect 3351 2023 3355 2031
rect 3359 2023 3363 2031
rect 1507 1993 1511 2001
rect 1520 1993 1524 2001
rect 1528 1993 1532 2001
rect 1536 1997 1540 2001
rect 1544 1993 1548 2001
rect 1557 1993 1561 2001
rect 1570 1993 1574 2001
rect 1578 1993 1582 2001
rect 1586 1993 1590 2001
rect 1594 1997 1598 2001
rect 1602 1993 1606 2001
rect 1615 1993 1619 2001
rect 1623 1993 1627 2001
rect 1631 1993 1635 2001
rect 1639 1993 1643 2001
rect 1652 1993 1656 2001
rect 1660 1993 1664 2001
rect 1668 1997 1672 2001
rect 1676 1993 1680 2001
rect 1689 1993 1693 2001
rect 1702 1993 1706 2001
rect 1710 1993 1714 2001
rect 1718 1993 1722 2001
rect 1726 1997 1730 2001
rect 1734 1993 1738 2001
rect 1747 1993 1751 2001
rect 1755 1993 1759 2001
rect 1763 1993 1767 2001
rect 1771 1993 1775 2001
rect 1784 1993 1788 2001
rect 1792 1993 1796 2001
rect 1800 1997 1804 2001
rect 1808 1993 1812 2001
rect 1821 1993 1825 2001
rect 1834 1993 1838 2001
rect 1842 1993 1846 2001
rect 1850 1993 1854 2001
rect 1858 1997 1862 2001
rect 1866 1993 1870 2001
rect 1879 1993 1883 2001
rect 1887 1993 1891 2001
rect 1895 1993 1899 2001
rect 2452 1993 2456 2001
rect 2465 1993 2469 2001
rect 2473 1993 2477 2001
rect 2481 1997 2485 2001
rect 2489 1993 2493 2001
rect 2502 1993 2506 2001
rect 2515 1993 2519 2001
rect 2523 1993 2527 2001
rect 2531 1993 2535 2001
rect 2539 1997 2543 2001
rect 2547 1993 2551 2001
rect 2560 1993 2564 2001
rect 2568 1993 2572 2001
rect 2576 1993 2580 2001
rect 2584 1993 2588 2001
rect 2597 1993 2601 2001
rect 2605 1993 2609 2001
rect 2613 1997 2617 2001
rect 2621 1993 2625 2001
rect 2634 1993 2638 2001
rect 2647 1993 2651 2001
rect 2655 1993 2659 2001
rect 2663 1993 2667 2001
rect 2671 1997 2675 2001
rect 2679 1993 2683 2001
rect 2692 1993 2696 2001
rect 2700 1993 2704 2001
rect 2708 1993 2712 2001
rect 2716 1993 2720 2001
rect 2729 1993 2733 2001
rect 2737 1993 2741 2001
rect 2745 1997 2749 2001
rect 2753 1993 2757 2001
rect 2766 1993 2770 2001
rect 2779 1993 2783 2001
rect 2787 1993 2791 2001
rect 2795 1993 2799 2001
rect 2803 1997 2807 2001
rect 2811 1993 2815 2001
rect 2824 1993 2828 2001
rect 2832 1993 2836 2001
rect 2840 1993 2844 2001
rect 1507 1853 1511 1861
rect 1520 1853 1524 1861
rect 1528 1853 1532 1861
rect 1536 1857 1540 1861
rect 1544 1853 1548 1861
rect 1557 1853 1561 1861
rect 1570 1853 1574 1861
rect 1578 1853 1582 1861
rect 1586 1853 1590 1861
rect 1594 1857 1598 1861
rect 1602 1853 1606 1861
rect 1615 1853 1619 1861
rect 1623 1853 1627 1861
rect 1631 1853 1635 1861
rect 1639 1853 1643 1861
rect 1652 1853 1656 1861
rect 1660 1853 1664 1861
rect 1668 1857 1672 1861
rect 1676 1853 1680 1861
rect 1689 1853 1693 1861
rect 1702 1853 1706 1861
rect 1710 1853 1714 1861
rect 1718 1853 1722 1861
rect 1726 1857 1730 1861
rect 1734 1853 1738 1861
rect 1747 1853 1751 1861
rect 1755 1853 1759 1861
rect 1763 1853 1767 1861
rect 1771 1853 1775 1861
rect 1784 1853 1788 1861
rect 1792 1853 1796 1861
rect 1800 1857 1804 1861
rect 1808 1853 1812 1861
rect 1821 1853 1825 1861
rect 1834 1853 1838 1861
rect 1842 1853 1846 1861
rect 1850 1853 1854 1861
rect 1858 1857 1862 1861
rect 1866 1853 1870 1861
rect 1879 1853 1883 1861
rect 1887 1853 1891 1861
rect 1895 1853 1899 1861
rect 2452 1853 2456 1861
rect 2465 1853 2469 1861
rect 2473 1853 2477 1861
rect 2481 1857 2485 1861
rect 2489 1853 2493 1861
rect 2502 1853 2506 1861
rect 2515 1853 2519 1861
rect 2523 1853 2527 1861
rect 2531 1853 2535 1861
rect 2539 1857 2543 1861
rect 2547 1853 2551 1861
rect 2560 1853 2564 1861
rect 2568 1853 2572 1861
rect 2576 1853 2580 1861
rect 2584 1853 2588 1861
rect 2597 1853 2601 1861
rect 2605 1853 2609 1861
rect 2613 1857 2617 1861
rect 2621 1853 2625 1861
rect 2634 1853 2638 1861
rect 2647 1853 2651 1861
rect 2655 1853 2659 1861
rect 2663 1853 2667 1861
rect 2671 1857 2675 1861
rect 2679 1853 2683 1861
rect 2692 1853 2696 1861
rect 2700 1853 2704 1861
rect 2708 1853 2712 1861
rect 2716 1853 2720 1861
rect 2729 1853 2733 1861
rect 2737 1853 2741 1861
rect 2745 1857 2749 1861
rect 2753 1853 2757 1861
rect 2766 1853 2770 1861
rect 2779 1853 2783 1861
rect 2787 1853 2791 1861
rect 2795 1853 2799 1861
rect 2803 1857 2807 1861
rect 2811 1853 2815 1861
rect 2824 1853 2828 1861
rect 2832 1853 2836 1861
rect 2840 1853 2844 1861
<< psubstratepcontact >>
rect 2689 4200 2693 4204
rect 2713 4200 2717 4204
rect 2767 4200 2771 4204
rect 2910 4200 2914 4204
rect 2667 4070 2671 4074
rect 2689 4070 2693 4074
rect 2713 4070 2717 4074
rect 2767 4070 2771 4074
rect 2816 4070 2820 4074
rect 2021 3699 2025 3703
rect 2049 3699 2053 3703
rect 2079 3699 2083 3703
rect 2153 3699 2157 3703
rect 2181 3699 2185 3703
rect 2211 3699 2215 3703
rect 2285 3699 2289 3703
rect 2313 3699 2317 3703
rect 2343 3699 2347 3703
rect 2417 3699 2421 3703
rect 2445 3699 2449 3703
rect 2475 3699 2479 3703
rect 2966 3699 2970 3703
rect 2994 3699 2998 3703
rect 3024 3699 3028 3703
rect 3098 3699 3102 3703
rect 3126 3699 3130 3703
rect 3156 3699 3160 3703
rect 3230 3699 3234 3703
rect 3258 3699 3262 3703
rect 3288 3699 3292 3703
rect 3362 3699 3366 3703
rect 3390 3699 3394 3703
rect 3420 3699 3424 3703
rect 1669 3666 1673 3670
rect 1697 3666 1701 3670
rect 1727 3666 1731 3670
rect 2614 3666 2618 3670
rect 2642 3666 2646 3670
rect 2672 3666 2676 3670
rect 2002 3613 2006 3617
rect 2037 3613 2041 3617
rect 2163 3613 2167 3617
rect 2187 3613 2191 3617
rect 2241 3613 2248 3617
rect 2268 3613 2272 3617
rect 2322 3613 2326 3617
rect 2947 3613 2951 3617
rect 2982 3613 2986 3617
rect 3108 3613 3112 3617
rect 3132 3613 3136 3617
rect 3186 3613 3193 3617
rect 3213 3613 3217 3617
rect 3267 3613 3271 3617
rect 1666 3564 1670 3568
rect 1696 3564 1700 3568
rect 1724 3564 1728 3568
rect 2611 3564 2615 3568
rect 2641 3564 2645 3568
rect 2669 3564 2673 3568
rect 2002 3481 2006 3485
rect 2037 3481 2041 3485
rect 2163 3481 2167 3485
rect 2187 3481 2191 3485
rect 2241 3481 2245 3485
rect 2268 3481 2272 3485
rect 2292 3481 2296 3485
rect 2947 3481 2951 3485
rect 2982 3481 2986 3485
rect 3108 3481 3112 3485
rect 3132 3481 3136 3485
rect 3186 3481 3190 3485
rect 3213 3481 3217 3485
rect 3237 3481 3241 3485
rect 2002 3349 2006 3353
rect 2037 3349 2041 3353
rect 2163 3349 2167 3353
rect 2187 3349 2191 3353
rect 2241 3349 2248 3353
rect 2268 3349 2272 3353
rect 2322 3349 2326 3353
rect 2358 3349 2362 3353
rect 2412 3349 2416 3353
rect 2947 3349 2951 3353
rect 2982 3349 2986 3353
rect 3108 3349 3112 3353
rect 3132 3349 3136 3353
rect 3186 3349 3193 3353
rect 3213 3349 3217 3353
rect 3267 3349 3271 3353
rect 3303 3349 3307 3353
rect 3357 3349 3361 3353
rect 2002 3217 2006 3221
rect 2037 3217 2041 3221
rect 2163 3217 2167 3221
rect 2187 3217 2191 3221
rect 2298 3217 2302 3221
rect 2947 3217 2951 3221
rect 2982 3217 2986 3221
rect 3108 3217 3112 3221
rect 3132 3217 3136 3221
rect 3243 3217 3247 3221
rect 1537 3164 1541 3168
rect 1565 3164 1569 3168
rect 1595 3164 1599 3168
rect 1669 3164 1673 3168
rect 1697 3164 1701 3168
rect 1727 3164 1731 3168
rect 1801 3164 1805 3168
rect 1829 3164 1833 3168
rect 1859 3164 1863 3168
rect 2482 3164 2486 3168
rect 2510 3164 2514 3168
rect 2540 3164 2544 3168
rect 2614 3164 2618 3168
rect 2642 3164 2646 3168
rect 2672 3164 2676 3168
rect 2746 3164 2750 3168
rect 2774 3164 2778 3168
rect 2804 3164 2808 3168
rect 2320 3052 2324 3056
rect 2348 3052 2352 3056
rect 2378 3052 2382 3056
rect 3265 3052 3269 3056
rect 3293 3052 3297 3056
rect 3323 3052 3327 3056
rect 1537 3022 1541 3026
rect 1565 3022 1569 3026
rect 1595 3022 1599 3026
rect 1669 3022 1673 3026
rect 1697 3022 1701 3026
rect 1727 3022 1731 3026
rect 1801 3022 1805 3026
rect 1829 3022 1833 3026
rect 1859 3022 1863 3026
rect 2482 3022 2486 3026
rect 2510 3022 2514 3026
rect 2540 3022 2544 3026
rect 2614 3022 2618 3026
rect 2642 3022 2646 3026
rect 2672 3022 2676 3026
rect 2746 3022 2750 3026
rect 2774 3022 2778 3026
rect 2804 3022 2808 3026
rect 2320 2966 2324 2970
rect 2348 2966 2352 2970
rect 2378 2966 2382 2970
rect 3265 2966 3269 2970
rect 3293 2966 3297 2970
rect 3323 2966 3327 2970
rect 1537 2936 1541 2940
rect 1565 2936 1569 2940
rect 1595 2936 1599 2940
rect 1669 2936 1673 2940
rect 1697 2936 1701 2940
rect 1727 2936 1731 2940
rect 1801 2936 1805 2940
rect 1829 2936 1833 2940
rect 1859 2936 1863 2940
rect 2482 2936 2486 2940
rect 2510 2936 2514 2940
rect 2540 2936 2544 2940
rect 2614 2936 2618 2940
rect 2642 2936 2646 2940
rect 2672 2936 2676 2940
rect 2746 2936 2750 2940
rect 2774 2936 2778 2940
rect 2804 2936 2808 2940
rect 1537 2796 1541 2800
rect 1565 2796 1569 2800
rect 1595 2796 1599 2800
rect 1669 2796 1673 2800
rect 1697 2796 1701 2800
rect 1727 2796 1731 2800
rect 1801 2796 1805 2800
rect 1829 2796 1833 2800
rect 1859 2796 1863 2800
rect 2482 2796 2486 2800
rect 2510 2796 2514 2800
rect 2540 2796 2544 2800
rect 2614 2796 2618 2800
rect 2642 2796 2646 2800
rect 2672 2796 2676 2800
rect 2746 2796 2750 2800
rect 2774 2796 2778 2800
rect 2804 2796 2808 2800
rect 2021 2717 2025 2721
rect 2049 2717 2053 2721
rect 2079 2717 2083 2721
rect 2153 2717 2157 2721
rect 2181 2717 2185 2721
rect 2211 2717 2215 2721
rect 2285 2717 2289 2721
rect 2313 2717 2317 2721
rect 2343 2717 2347 2721
rect 2417 2717 2421 2721
rect 2445 2717 2449 2721
rect 2475 2717 2479 2721
rect 2966 2717 2970 2721
rect 2994 2717 2998 2721
rect 3024 2717 3028 2721
rect 3098 2717 3102 2721
rect 3126 2717 3130 2721
rect 3156 2717 3160 2721
rect 3230 2717 3234 2721
rect 3258 2717 3262 2721
rect 3288 2717 3292 2721
rect 3362 2717 3366 2721
rect 3390 2717 3394 2721
rect 3420 2717 3424 2721
rect 1669 2684 1673 2688
rect 1697 2684 1701 2688
rect 1727 2684 1731 2688
rect 2614 2684 2618 2688
rect 2642 2684 2646 2688
rect 2672 2684 2676 2688
rect 2002 2631 2006 2635
rect 2037 2631 2041 2635
rect 2163 2631 2167 2635
rect 2187 2631 2191 2635
rect 2241 2631 2248 2635
rect 2268 2631 2272 2635
rect 2322 2631 2326 2635
rect 2947 2631 2951 2635
rect 2982 2631 2986 2635
rect 3108 2631 3112 2635
rect 3132 2631 3136 2635
rect 3186 2631 3193 2635
rect 3213 2631 3217 2635
rect 3267 2631 3271 2635
rect 1666 2582 1670 2586
rect 1696 2582 1700 2586
rect 1724 2582 1728 2586
rect 2611 2582 2615 2586
rect 2641 2582 2645 2586
rect 2669 2582 2673 2586
rect 2002 2499 2006 2503
rect 2037 2499 2041 2503
rect 2163 2499 2167 2503
rect 2187 2499 2191 2503
rect 2241 2499 2245 2503
rect 2268 2499 2272 2503
rect 2292 2499 2296 2503
rect 2947 2499 2951 2503
rect 2982 2499 2986 2503
rect 3108 2499 3112 2503
rect 3132 2499 3136 2503
rect 3186 2499 3190 2503
rect 3213 2499 3217 2503
rect 3237 2499 3241 2503
rect 2002 2367 2006 2371
rect 2037 2367 2041 2371
rect 2163 2367 2167 2371
rect 2187 2367 2191 2371
rect 2241 2367 2248 2371
rect 2268 2367 2272 2371
rect 2322 2367 2326 2371
rect 2358 2367 2362 2371
rect 2412 2367 2416 2371
rect 2947 2367 2951 2371
rect 2982 2367 2986 2371
rect 3108 2367 3112 2371
rect 3132 2367 3136 2371
rect 3186 2367 3193 2371
rect 3213 2367 3217 2371
rect 3267 2367 3271 2371
rect 3303 2367 3307 2371
rect 3357 2367 3361 2371
rect 2002 2235 2006 2239
rect 2037 2235 2041 2239
rect 2163 2235 2167 2239
rect 2187 2235 2191 2239
rect 2298 2235 2302 2239
rect 2947 2235 2951 2239
rect 2982 2235 2986 2239
rect 3108 2235 3112 2239
rect 3132 2235 3136 2239
rect 3243 2235 3247 2239
rect 1537 2182 1541 2186
rect 1565 2182 1569 2186
rect 1595 2182 1599 2186
rect 1669 2182 1673 2186
rect 1697 2182 1701 2186
rect 1727 2182 1731 2186
rect 1801 2182 1805 2186
rect 1829 2182 1833 2186
rect 1859 2182 1863 2186
rect 2482 2182 2486 2186
rect 2510 2182 2514 2186
rect 2540 2182 2544 2186
rect 2614 2182 2618 2186
rect 2642 2182 2646 2186
rect 2672 2182 2676 2186
rect 2746 2182 2750 2186
rect 2774 2182 2778 2186
rect 2804 2182 2808 2186
rect 2320 2070 2324 2074
rect 2348 2070 2352 2074
rect 2378 2070 2382 2074
rect 3265 2070 3269 2074
rect 3293 2070 3297 2074
rect 3323 2070 3327 2074
rect 1537 2040 1541 2044
rect 1565 2040 1569 2044
rect 1595 2040 1599 2044
rect 1669 2040 1673 2044
rect 1697 2040 1701 2044
rect 1727 2040 1731 2044
rect 1801 2040 1805 2044
rect 1829 2040 1833 2044
rect 1859 2040 1863 2044
rect 2482 2040 2486 2044
rect 2510 2040 2514 2044
rect 2540 2040 2544 2044
rect 2614 2040 2618 2044
rect 2642 2040 2646 2044
rect 2672 2040 2676 2044
rect 2746 2040 2750 2044
rect 2774 2040 2778 2044
rect 2804 2040 2808 2044
rect 2320 1984 2324 1988
rect 2348 1984 2352 1988
rect 2378 1984 2382 1988
rect 3265 1984 3269 1988
rect 3293 1984 3297 1988
rect 3323 1984 3327 1988
rect 1537 1954 1541 1958
rect 1565 1954 1569 1958
rect 1595 1954 1599 1958
rect 1669 1954 1673 1958
rect 1697 1954 1701 1958
rect 1727 1954 1731 1958
rect 1801 1954 1805 1958
rect 1829 1954 1833 1958
rect 1859 1954 1863 1958
rect 2482 1954 2486 1958
rect 2510 1954 2514 1958
rect 2540 1954 2544 1958
rect 2614 1954 2618 1958
rect 2642 1954 2646 1958
rect 2672 1954 2676 1958
rect 2746 1954 2750 1958
rect 2774 1954 2778 1958
rect 2804 1954 2808 1958
rect 1537 1814 1541 1818
rect 1565 1814 1569 1818
rect 1595 1814 1599 1818
rect 1669 1814 1673 1818
rect 1697 1814 1701 1818
rect 1727 1814 1731 1818
rect 1801 1814 1805 1818
rect 1829 1814 1833 1818
rect 1859 1814 1863 1818
rect 2482 1814 2486 1818
rect 2510 1814 2514 1818
rect 2540 1814 2544 1818
rect 2614 1814 2618 1818
rect 2642 1814 2646 1818
rect 2672 1814 2676 1818
rect 2746 1814 2750 1818
rect 2774 1814 2778 1818
rect 2804 1814 2808 1818
<< nsubstratencontact >>
rect 2689 4280 2693 4284
rect 2713 4280 2717 4284
rect 2767 4280 2771 4284
rect 2910 4280 2914 4284
rect 2667 4150 2671 4154
rect 2689 4150 2693 4154
rect 2713 4150 2717 4154
rect 2767 4150 2771 4154
rect 2816 4150 2820 4154
rect 2713 4020 2717 4024
rect 2021 3756 2025 3760
rect 2049 3756 2053 3760
rect 2079 3756 2083 3760
rect 2116 3756 2120 3760
rect 2153 3756 2157 3760
rect 2181 3756 2185 3760
rect 2211 3756 2215 3760
rect 2248 3756 2252 3760
rect 2285 3756 2289 3760
rect 2313 3756 2317 3760
rect 2343 3756 2347 3760
rect 2380 3756 2384 3760
rect 2417 3756 2421 3760
rect 2445 3756 2449 3760
rect 2475 3756 2479 3760
rect 2512 3756 2516 3760
rect 2966 3756 2970 3760
rect 2994 3756 2998 3760
rect 3024 3756 3028 3760
rect 3061 3756 3065 3760
rect 3098 3756 3102 3760
rect 3126 3756 3130 3760
rect 3156 3756 3160 3760
rect 3193 3756 3197 3760
rect 3230 3756 3234 3760
rect 3258 3756 3262 3760
rect 3288 3756 3292 3760
rect 3325 3756 3329 3760
rect 3362 3756 3366 3760
rect 3390 3756 3394 3760
rect 3420 3756 3424 3760
rect 3457 3756 3461 3760
rect 1669 3723 1673 3727
rect 1697 3723 1701 3727
rect 1727 3723 1731 3727
rect 1764 3723 1768 3727
rect 2614 3723 2618 3727
rect 2642 3723 2646 3727
rect 2672 3723 2676 3727
rect 2709 3723 2713 3727
rect 2011 3679 2015 3683
rect 2040 3679 2044 3683
rect 2065 3679 2069 3683
rect 2107 3679 2111 3683
rect 2163 3679 2167 3683
rect 2187 3679 2191 3683
rect 2241 3679 2245 3683
rect 2268 3679 2272 3683
rect 2322 3679 2326 3683
rect 2956 3679 2960 3683
rect 2985 3679 2989 3683
rect 3010 3679 3014 3683
rect 3052 3679 3056 3683
rect 3108 3679 3112 3683
rect 3132 3679 3136 3683
rect 3186 3679 3190 3683
rect 3213 3679 3217 3683
rect 3267 3679 3271 3683
rect 1629 3621 1633 3625
rect 1666 3621 1670 3625
rect 1696 3621 1700 3625
rect 1724 3621 1728 3625
rect 2574 3621 2578 3625
rect 2611 3621 2615 3625
rect 2641 3621 2645 3625
rect 2669 3621 2673 3625
rect 2011 3547 2015 3551
rect 2040 3547 2044 3551
rect 2065 3547 2069 3551
rect 2107 3547 2111 3551
rect 2163 3547 2167 3551
rect 2187 3547 2191 3551
rect 2241 3547 2245 3551
rect 2268 3547 2272 3551
rect 2330 3547 2334 3551
rect 2956 3547 2960 3551
rect 2985 3547 2989 3551
rect 3010 3547 3014 3551
rect 3052 3547 3056 3551
rect 3108 3547 3112 3551
rect 3132 3547 3136 3551
rect 3186 3547 3190 3551
rect 3213 3547 3217 3551
rect 3275 3547 3279 3551
rect 2011 3415 2015 3419
rect 2040 3415 2044 3419
rect 2065 3415 2069 3419
rect 2107 3415 2111 3419
rect 2163 3415 2167 3419
rect 2187 3415 2191 3419
rect 2241 3415 2245 3419
rect 2268 3415 2272 3419
rect 2322 3415 2326 3419
rect 2330 3415 2334 3419
rect 2358 3415 2362 3419
rect 2412 3415 2416 3419
rect 2956 3415 2960 3419
rect 2985 3415 2989 3419
rect 3010 3415 3014 3419
rect 3052 3415 3056 3419
rect 3108 3415 3112 3419
rect 3132 3415 3136 3419
rect 3186 3415 3190 3419
rect 3213 3415 3217 3419
rect 3267 3415 3271 3419
rect 3275 3415 3279 3419
rect 3303 3415 3307 3419
rect 3357 3415 3361 3419
rect 2011 3283 2015 3287
rect 2040 3283 2044 3287
rect 2065 3283 2069 3287
rect 2107 3283 2111 3287
rect 2163 3283 2167 3287
rect 2187 3283 2191 3287
rect 2241 3283 2245 3287
rect 2268 3283 2272 3287
rect 2358 3283 2362 3287
rect 2956 3283 2960 3287
rect 2985 3283 2989 3287
rect 3010 3283 3014 3287
rect 3052 3283 3056 3287
rect 3108 3283 3112 3287
rect 3132 3283 3136 3287
rect 3186 3283 3190 3287
rect 3213 3283 3217 3287
rect 3303 3283 3307 3287
rect 1537 3221 1541 3225
rect 1565 3221 1569 3225
rect 1595 3221 1599 3225
rect 1632 3221 1636 3225
rect 1669 3221 1673 3225
rect 1697 3221 1701 3225
rect 1727 3221 1731 3225
rect 1764 3221 1768 3225
rect 1801 3221 1805 3225
rect 1829 3221 1833 3225
rect 1859 3221 1863 3225
rect 1896 3221 1900 3225
rect 2482 3221 2486 3225
rect 2510 3221 2514 3225
rect 2540 3221 2544 3225
rect 2577 3221 2581 3225
rect 2614 3221 2618 3225
rect 2642 3221 2646 3225
rect 2672 3221 2676 3225
rect 2709 3221 2713 3225
rect 2746 3221 2750 3225
rect 2774 3221 2778 3225
rect 2804 3221 2808 3225
rect 2841 3221 2845 3225
rect 2011 3151 2015 3155
rect 2040 3151 2044 3155
rect 2065 3151 2069 3155
rect 2107 3151 2111 3155
rect 2187 3151 2191 3155
rect 2241 3151 2245 3155
rect 2272 3151 2276 3155
rect 2301 3151 2305 3155
rect 2326 3151 2330 3155
rect 2368 3151 2372 3155
rect 2956 3151 2960 3155
rect 2985 3151 2989 3155
rect 3010 3151 3014 3155
rect 3052 3151 3056 3155
rect 3132 3151 3136 3155
rect 3186 3151 3190 3155
rect 3217 3151 3221 3155
rect 3246 3151 3250 3155
rect 3271 3151 3275 3155
rect 3313 3151 3317 3155
rect 2320 3109 2324 3113
rect 2348 3109 2352 3113
rect 2378 3109 2382 3113
rect 2415 3109 2419 3113
rect 3265 3109 3269 3113
rect 3293 3109 3297 3113
rect 3323 3109 3327 3113
rect 3360 3109 3364 3113
rect 1537 3079 1541 3083
rect 1565 3079 1569 3083
rect 1595 3079 1599 3083
rect 1632 3079 1636 3083
rect 1669 3079 1673 3083
rect 1697 3079 1701 3083
rect 1727 3079 1731 3083
rect 1764 3079 1768 3083
rect 1801 3079 1805 3083
rect 1829 3079 1833 3083
rect 1859 3079 1863 3083
rect 1896 3079 1900 3083
rect 2482 3079 2486 3083
rect 2510 3079 2514 3083
rect 2540 3079 2544 3083
rect 2577 3079 2581 3083
rect 2614 3079 2618 3083
rect 2642 3079 2646 3083
rect 2672 3079 2676 3083
rect 2709 3079 2713 3083
rect 2746 3079 2750 3083
rect 2774 3079 2778 3083
rect 2804 3079 2808 3083
rect 2841 3079 2845 3083
rect 2320 3023 2324 3027
rect 2348 3023 2352 3027
rect 2378 3023 2382 3027
rect 2415 3023 2419 3027
rect 3265 3023 3269 3027
rect 3293 3023 3297 3027
rect 3323 3023 3327 3027
rect 3360 3023 3364 3027
rect 1537 2993 1541 2997
rect 1565 2993 1569 2997
rect 1595 2993 1599 2997
rect 1632 2993 1636 2997
rect 1669 2993 1673 2997
rect 1697 2993 1701 2997
rect 1727 2993 1731 2997
rect 1764 2993 1768 2997
rect 1801 2993 1805 2997
rect 1829 2993 1833 2997
rect 1859 2993 1863 2997
rect 1896 2993 1900 2997
rect 2482 2993 2486 2997
rect 2510 2993 2514 2997
rect 2540 2993 2544 2997
rect 2577 2993 2581 2997
rect 2614 2993 2618 2997
rect 2642 2993 2646 2997
rect 2672 2993 2676 2997
rect 2709 2993 2713 2997
rect 2746 2993 2750 2997
rect 2774 2993 2778 2997
rect 2804 2993 2808 2997
rect 2841 2993 2845 2997
rect 1537 2853 1541 2857
rect 1565 2853 1569 2857
rect 1595 2853 1599 2857
rect 1632 2853 1636 2857
rect 1669 2853 1673 2857
rect 1697 2853 1701 2857
rect 1727 2853 1731 2857
rect 1764 2853 1768 2857
rect 1801 2853 1805 2857
rect 1829 2853 1833 2857
rect 1859 2853 1863 2857
rect 1896 2853 1900 2857
rect 2482 2853 2486 2857
rect 2510 2853 2514 2857
rect 2540 2853 2544 2857
rect 2577 2853 2581 2857
rect 2614 2853 2618 2857
rect 2642 2853 2646 2857
rect 2672 2853 2676 2857
rect 2709 2853 2713 2857
rect 2746 2853 2750 2857
rect 2774 2853 2778 2857
rect 2804 2853 2808 2857
rect 2841 2853 2845 2857
rect 2021 2774 2025 2778
rect 2049 2774 2053 2778
rect 2079 2774 2083 2778
rect 2116 2774 2120 2778
rect 2153 2774 2157 2778
rect 2181 2774 2185 2778
rect 2211 2774 2215 2778
rect 2248 2774 2252 2778
rect 2285 2774 2289 2778
rect 2313 2774 2317 2778
rect 2343 2774 2347 2778
rect 2380 2774 2384 2778
rect 2417 2774 2421 2778
rect 2445 2774 2449 2778
rect 2475 2774 2479 2778
rect 2512 2774 2516 2778
rect 2966 2774 2970 2778
rect 2994 2774 2998 2778
rect 3024 2774 3028 2778
rect 3061 2774 3065 2778
rect 3098 2774 3102 2778
rect 3126 2774 3130 2778
rect 3156 2774 3160 2778
rect 3193 2774 3197 2778
rect 3230 2774 3234 2778
rect 3258 2774 3262 2778
rect 3288 2774 3292 2778
rect 3325 2774 3329 2778
rect 3362 2774 3366 2778
rect 3390 2774 3394 2778
rect 3420 2774 3424 2778
rect 3457 2774 3461 2778
rect 1669 2741 1673 2745
rect 1697 2741 1701 2745
rect 1727 2741 1731 2745
rect 1764 2741 1768 2745
rect 2614 2741 2618 2745
rect 2642 2741 2646 2745
rect 2672 2741 2676 2745
rect 2709 2741 2713 2745
rect 2011 2697 2015 2701
rect 2040 2697 2044 2701
rect 2065 2697 2069 2701
rect 2107 2697 2111 2701
rect 2163 2697 2167 2701
rect 2187 2697 2191 2701
rect 2241 2697 2245 2701
rect 2268 2697 2272 2701
rect 2322 2697 2326 2701
rect 2956 2697 2960 2701
rect 2985 2697 2989 2701
rect 3010 2697 3014 2701
rect 3052 2697 3056 2701
rect 3108 2697 3112 2701
rect 3132 2697 3136 2701
rect 3186 2697 3190 2701
rect 3213 2697 3217 2701
rect 3267 2697 3271 2701
rect 1629 2639 1633 2643
rect 1666 2639 1670 2643
rect 1696 2639 1700 2643
rect 1724 2639 1728 2643
rect 2574 2639 2578 2643
rect 2611 2639 2615 2643
rect 2641 2639 2645 2643
rect 2669 2639 2673 2643
rect 2011 2565 2015 2569
rect 2040 2565 2044 2569
rect 2065 2565 2069 2569
rect 2107 2565 2111 2569
rect 2163 2565 2167 2569
rect 2187 2565 2191 2569
rect 2241 2565 2245 2569
rect 2268 2565 2272 2569
rect 2330 2565 2334 2569
rect 2956 2565 2960 2569
rect 2985 2565 2989 2569
rect 3010 2565 3014 2569
rect 3052 2565 3056 2569
rect 3108 2565 3112 2569
rect 3132 2565 3136 2569
rect 3186 2565 3190 2569
rect 3213 2565 3217 2569
rect 3275 2565 3279 2569
rect 2011 2433 2015 2437
rect 2040 2433 2044 2437
rect 2065 2433 2069 2437
rect 2107 2433 2111 2437
rect 2163 2433 2167 2437
rect 2187 2433 2191 2437
rect 2241 2433 2245 2437
rect 2268 2433 2272 2437
rect 2322 2433 2326 2437
rect 2330 2433 2334 2437
rect 2358 2433 2362 2437
rect 2412 2433 2416 2437
rect 2956 2433 2960 2437
rect 2985 2433 2989 2437
rect 3010 2433 3014 2437
rect 3052 2433 3056 2437
rect 3108 2433 3112 2437
rect 3132 2433 3136 2437
rect 3186 2433 3190 2437
rect 3213 2433 3217 2437
rect 3267 2433 3271 2437
rect 3275 2433 3279 2437
rect 3303 2433 3307 2437
rect 3357 2433 3361 2437
rect 2011 2301 2015 2305
rect 2040 2301 2044 2305
rect 2065 2301 2069 2305
rect 2107 2301 2111 2305
rect 2163 2301 2167 2305
rect 2187 2301 2191 2305
rect 2241 2301 2245 2305
rect 2268 2301 2272 2305
rect 2358 2301 2362 2305
rect 2956 2301 2960 2305
rect 2985 2301 2989 2305
rect 3010 2301 3014 2305
rect 3052 2301 3056 2305
rect 3108 2301 3112 2305
rect 3132 2301 3136 2305
rect 3186 2301 3190 2305
rect 3213 2301 3217 2305
rect 3303 2301 3307 2305
rect 1537 2239 1541 2243
rect 1565 2239 1569 2243
rect 1595 2239 1599 2243
rect 1632 2239 1636 2243
rect 1669 2239 1673 2243
rect 1697 2239 1701 2243
rect 1727 2239 1731 2243
rect 1764 2239 1768 2243
rect 1801 2239 1805 2243
rect 1829 2239 1833 2243
rect 1859 2239 1863 2243
rect 1896 2239 1900 2243
rect 2482 2239 2486 2243
rect 2510 2239 2514 2243
rect 2540 2239 2544 2243
rect 2577 2239 2581 2243
rect 2614 2239 2618 2243
rect 2642 2239 2646 2243
rect 2672 2239 2676 2243
rect 2709 2239 2713 2243
rect 2746 2239 2750 2243
rect 2774 2239 2778 2243
rect 2804 2239 2808 2243
rect 2841 2239 2845 2243
rect 2011 2169 2015 2173
rect 2040 2169 2044 2173
rect 2065 2169 2069 2173
rect 2107 2169 2111 2173
rect 2187 2169 2191 2173
rect 2241 2169 2245 2173
rect 2272 2169 2276 2173
rect 2301 2169 2305 2173
rect 2326 2169 2330 2173
rect 2368 2169 2372 2173
rect 2956 2169 2960 2173
rect 2985 2169 2989 2173
rect 3010 2169 3014 2173
rect 3052 2169 3056 2173
rect 3132 2169 3136 2173
rect 3186 2169 3190 2173
rect 3217 2169 3221 2173
rect 3246 2169 3250 2173
rect 3271 2169 3275 2173
rect 3313 2169 3317 2173
rect 2320 2127 2324 2131
rect 2348 2127 2352 2131
rect 2378 2127 2382 2131
rect 2415 2127 2419 2131
rect 3265 2127 3269 2131
rect 3293 2127 3297 2131
rect 3323 2127 3327 2131
rect 3360 2127 3364 2131
rect 1537 2097 1541 2101
rect 1565 2097 1569 2101
rect 1595 2097 1599 2101
rect 1632 2097 1636 2101
rect 1669 2097 1673 2101
rect 1697 2097 1701 2101
rect 1727 2097 1731 2101
rect 1764 2097 1768 2101
rect 1801 2097 1805 2101
rect 1829 2097 1833 2101
rect 1859 2097 1863 2101
rect 1896 2097 1900 2101
rect 2482 2097 2486 2101
rect 2510 2097 2514 2101
rect 2540 2097 2544 2101
rect 2577 2097 2581 2101
rect 2614 2097 2618 2101
rect 2642 2097 2646 2101
rect 2672 2097 2676 2101
rect 2709 2097 2713 2101
rect 2746 2097 2750 2101
rect 2774 2097 2778 2101
rect 2804 2097 2808 2101
rect 2841 2097 2845 2101
rect 2320 2041 2324 2045
rect 2348 2041 2352 2045
rect 2378 2041 2382 2045
rect 2415 2041 2419 2045
rect 3265 2041 3269 2045
rect 3293 2041 3297 2045
rect 3323 2041 3327 2045
rect 3360 2041 3364 2045
rect 1537 2011 1541 2015
rect 1565 2011 1569 2015
rect 1595 2011 1599 2015
rect 1632 2011 1636 2015
rect 1669 2011 1673 2015
rect 1697 2011 1701 2015
rect 1727 2011 1731 2015
rect 1764 2011 1768 2015
rect 1801 2011 1805 2015
rect 1829 2011 1833 2015
rect 1859 2011 1863 2015
rect 1896 2011 1900 2015
rect 2482 2011 2486 2015
rect 2510 2011 2514 2015
rect 2540 2011 2544 2015
rect 2577 2011 2581 2015
rect 2614 2011 2618 2015
rect 2642 2011 2646 2015
rect 2672 2011 2676 2015
rect 2709 2011 2713 2015
rect 2746 2011 2750 2015
rect 2774 2011 2778 2015
rect 2804 2011 2808 2015
rect 2841 2011 2845 2015
rect 1537 1871 1541 1875
rect 1565 1871 1569 1875
rect 1595 1871 1599 1875
rect 1632 1871 1636 1875
rect 1669 1871 1673 1875
rect 1697 1871 1701 1875
rect 1727 1871 1731 1875
rect 1764 1871 1768 1875
rect 1801 1871 1805 1875
rect 1829 1871 1833 1875
rect 1859 1871 1863 1875
rect 1896 1871 1900 1875
rect 2482 1871 2486 1875
rect 2510 1871 2514 1875
rect 2540 1871 2544 1875
rect 2577 1871 2581 1875
rect 2614 1871 2618 1875
rect 2642 1871 2646 1875
rect 2672 1871 2676 1875
rect 2709 1871 2713 1875
rect 2746 1871 2750 1875
rect 2774 1871 2778 1875
rect 2804 1871 2808 1875
rect 2841 1871 2845 1875
<< polysilicon >>
rect 2701 4276 2703 4278
rect 2727 4270 2729 4274
rect 2755 4276 2757 4278
rect 2732 4270 2734 4273
rect 2701 4254 2703 4268
rect 2887 4273 2889 4276
rect 2940 4273 2942 4276
rect 2727 4259 2729 4262
rect 2732 4260 2734 4262
rect 2728 4255 2729 4259
rect 2727 4250 2729 4255
rect 2732 4250 2734 4252
rect 2701 4248 2703 4250
rect 2755 4246 2757 4268
rect 2727 4244 2729 4246
rect 2732 4241 2734 4246
rect 2755 4240 2757 4242
rect 2887 4235 2889 4243
rect 2940 4235 2942 4243
rect 2887 4223 2889 4231
rect 2940 4223 2942 4231
rect 2887 4209 2889 4211
rect 2940 4209 2942 4211
rect 2727 4190 2729 4193
rect 2732 4190 2734 4193
rect 2727 4174 2729 4186
rect 2732 4184 2734 4186
rect 2732 4174 2734 4176
rect 2727 4164 2729 4166
rect 2732 4161 2734 4166
rect 2679 4146 2681 4148
rect 2701 4146 2703 4148
rect 2727 4140 2729 4144
rect 2755 4146 2757 4148
rect 2732 4140 2734 4143
rect 2679 4124 2681 4138
rect 2701 4124 2703 4138
rect 2793 4143 2795 4146
rect 2846 4143 2848 4146
rect 2727 4129 2729 4132
rect 2732 4130 2734 4132
rect 2728 4125 2729 4129
rect 2727 4120 2729 4125
rect 2732 4120 2734 4122
rect 2679 4118 2681 4120
rect 2701 4118 2703 4120
rect 2755 4116 2757 4138
rect 2727 4114 2729 4116
rect 2732 4111 2734 4116
rect 2755 4110 2757 4112
rect 2793 4105 2795 4113
rect 2846 4105 2848 4113
rect 2793 4093 2795 4101
rect 2846 4093 2848 4101
rect 2793 4079 2795 4081
rect 2846 4079 2848 4081
rect 2727 4060 2729 4063
rect 2732 4060 2734 4063
rect 2727 4044 2729 4056
rect 2732 4054 2734 4056
rect 2732 4044 2734 4046
rect 2727 4034 2729 4036
rect 2732 4031 2734 4036
rect 1996 3746 1998 3748
rect 2001 3746 2003 3749
rect 2017 3746 2019 3748
rect 2033 3746 2035 3748
rect 2038 3746 2040 3749
rect 2059 3746 2061 3749
rect 2075 3746 2077 3749
rect 2091 3746 2093 3748
rect 2096 3746 2098 3749
rect 2112 3746 2114 3748
rect 2128 3746 2130 3748
rect 2133 3746 2135 3749
rect 2149 3746 2151 3748
rect 2165 3746 2167 3748
rect 2170 3746 2172 3749
rect 2191 3746 2193 3749
rect 2207 3746 2209 3749
rect 2223 3746 2225 3748
rect 2228 3746 2230 3749
rect 2244 3746 2246 3748
rect 2260 3746 2262 3748
rect 2265 3746 2267 3749
rect 2281 3746 2283 3748
rect 2297 3746 2299 3748
rect 2302 3746 2304 3749
rect 2323 3746 2325 3749
rect 2339 3746 2341 3749
rect 2355 3746 2357 3748
rect 2360 3746 2362 3749
rect 2376 3746 2378 3748
rect 2392 3746 2394 3748
rect 2397 3746 2399 3749
rect 2413 3746 2415 3748
rect 2429 3746 2431 3748
rect 2434 3746 2436 3749
rect 2455 3746 2457 3749
rect 2471 3746 2473 3749
rect 2487 3746 2489 3748
rect 2492 3746 2494 3749
rect 2508 3746 2510 3748
rect 2941 3746 2943 3748
rect 2946 3746 2948 3749
rect 2962 3746 2964 3748
rect 2978 3746 2980 3748
rect 2983 3746 2985 3749
rect 3004 3746 3006 3749
rect 3020 3746 3022 3749
rect 3036 3746 3038 3748
rect 3041 3746 3043 3749
rect 3057 3746 3059 3748
rect 3073 3746 3075 3748
rect 3078 3746 3080 3749
rect 3094 3746 3096 3748
rect 3110 3746 3112 3748
rect 3115 3746 3117 3749
rect 3136 3746 3138 3749
rect 3152 3746 3154 3749
rect 3168 3746 3170 3748
rect 3173 3746 3175 3749
rect 3189 3746 3191 3748
rect 3205 3746 3207 3748
rect 3210 3746 3212 3749
rect 3226 3746 3228 3748
rect 3242 3746 3244 3748
rect 3247 3746 3249 3749
rect 3268 3746 3270 3749
rect 3284 3746 3286 3749
rect 3300 3746 3302 3748
rect 3305 3746 3307 3749
rect 3321 3746 3323 3748
rect 3337 3746 3339 3748
rect 3342 3746 3344 3749
rect 3358 3746 3360 3748
rect 3374 3746 3376 3748
rect 3379 3746 3381 3749
rect 3400 3746 3402 3749
rect 3416 3746 3418 3749
rect 3432 3746 3434 3748
rect 3437 3746 3439 3749
rect 3453 3746 3455 3748
rect 1996 3733 1998 3738
rect 2001 3736 2003 3738
rect 1996 3719 1998 3729
rect 2001 3719 2003 3726
rect 2017 3719 2019 3738
rect 2033 3729 2035 3738
rect 2038 3736 2040 3738
rect 2059 3736 2061 3738
rect 2075 3735 2077 3738
rect 2033 3719 2035 3722
rect 2038 3719 2040 3721
rect 2059 3719 2061 3721
rect 2075 3719 2077 3731
rect 2091 3729 2093 3738
rect 2096 3736 2098 3738
rect 2112 3730 2114 3738
rect 2128 3733 2130 3738
rect 2133 3736 2135 3738
rect 2091 3719 2093 3722
rect 2096 3719 2098 3721
rect 2112 3719 2114 3726
rect 2128 3719 2130 3729
rect 2133 3719 2135 3726
rect 2149 3719 2151 3738
rect 2165 3729 2167 3738
rect 2170 3736 2172 3738
rect 2191 3736 2193 3738
rect 2207 3735 2209 3738
rect 2165 3719 2167 3722
rect 2170 3719 2172 3721
rect 2191 3719 2193 3721
rect 2207 3719 2209 3731
rect 2223 3729 2225 3738
rect 2228 3736 2230 3738
rect 2244 3730 2246 3738
rect 2260 3733 2262 3738
rect 2265 3736 2267 3738
rect 2223 3719 2225 3722
rect 2228 3719 2230 3721
rect 2244 3719 2246 3726
rect 2260 3719 2262 3729
rect 2265 3719 2267 3726
rect 2281 3719 2283 3738
rect 2297 3729 2299 3738
rect 2302 3736 2304 3738
rect 2323 3736 2325 3738
rect 2339 3735 2341 3738
rect 2297 3719 2299 3722
rect 2302 3719 2304 3721
rect 2323 3719 2325 3721
rect 2339 3719 2341 3731
rect 2355 3729 2357 3738
rect 2360 3736 2362 3738
rect 2376 3730 2378 3738
rect 2392 3733 2394 3738
rect 2397 3736 2399 3738
rect 2355 3719 2357 3722
rect 2360 3719 2362 3721
rect 2376 3719 2378 3726
rect 2392 3719 2394 3729
rect 2397 3719 2399 3726
rect 2413 3719 2415 3738
rect 2429 3729 2431 3738
rect 2434 3736 2436 3738
rect 2455 3736 2457 3738
rect 2471 3735 2473 3738
rect 2429 3719 2431 3722
rect 2434 3719 2436 3721
rect 2455 3719 2457 3721
rect 2471 3719 2473 3731
rect 2487 3729 2489 3738
rect 2492 3736 2494 3738
rect 2508 3730 2510 3738
rect 2941 3733 2943 3738
rect 2946 3736 2948 3738
rect 2487 3719 2489 3722
rect 2492 3719 2494 3721
rect 2508 3719 2510 3726
rect 1644 3713 1646 3715
rect 1649 3713 1651 3716
rect 1665 3713 1667 3715
rect 1681 3713 1683 3715
rect 1686 3713 1688 3716
rect 1707 3713 1709 3716
rect 1723 3713 1725 3716
rect 1739 3713 1741 3715
rect 1744 3713 1746 3716
rect 2941 3719 2943 3729
rect 2946 3719 2948 3726
rect 2962 3719 2964 3738
rect 2978 3729 2980 3738
rect 2983 3736 2985 3738
rect 3004 3736 3006 3738
rect 3020 3735 3022 3738
rect 2978 3719 2980 3722
rect 2983 3719 2985 3721
rect 3004 3719 3006 3721
rect 3020 3719 3022 3731
rect 3036 3729 3038 3738
rect 3041 3736 3043 3738
rect 3057 3730 3059 3738
rect 3073 3733 3075 3738
rect 3078 3736 3080 3738
rect 3036 3719 3038 3722
rect 3041 3719 3043 3721
rect 3057 3719 3059 3726
rect 3073 3719 3075 3729
rect 3078 3719 3080 3726
rect 3094 3719 3096 3738
rect 3110 3729 3112 3738
rect 3115 3736 3117 3738
rect 3136 3736 3138 3738
rect 3152 3735 3154 3738
rect 3110 3719 3112 3722
rect 3115 3719 3117 3721
rect 3136 3719 3138 3721
rect 3152 3719 3154 3731
rect 3168 3729 3170 3738
rect 3173 3736 3175 3738
rect 3189 3730 3191 3738
rect 3205 3733 3207 3738
rect 3210 3736 3212 3738
rect 3168 3719 3170 3722
rect 3173 3719 3175 3721
rect 3189 3719 3191 3726
rect 3205 3719 3207 3729
rect 3210 3719 3212 3726
rect 3226 3719 3228 3738
rect 3242 3729 3244 3738
rect 3247 3736 3249 3738
rect 3268 3736 3270 3738
rect 3284 3735 3286 3738
rect 3242 3719 3244 3722
rect 3247 3719 3249 3721
rect 3268 3719 3270 3721
rect 3284 3719 3286 3731
rect 3300 3729 3302 3738
rect 3305 3736 3307 3738
rect 3321 3730 3323 3738
rect 3337 3733 3339 3738
rect 3342 3736 3344 3738
rect 3300 3719 3302 3722
rect 3305 3719 3307 3721
rect 3321 3719 3323 3726
rect 3337 3719 3339 3729
rect 3342 3719 3344 3726
rect 3358 3719 3360 3738
rect 3374 3729 3376 3738
rect 3379 3736 3381 3738
rect 3400 3736 3402 3738
rect 3416 3735 3418 3738
rect 3374 3719 3376 3722
rect 3379 3719 3381 3721
rect 3400 3719 3402 3721
rect 3416 3719 3418 3731
rect 3432 3729 3434 3738
rect 3437 3736 3439 3738
rect 3453 3730 3455 3738
rect 3432 3719 3434 3722
rect 3437 3719 3439 3721
rect 3453 3719 3455 3726
rect 1760 3713 1762 3715
rect 1996 3713 1998 3715
rect 2001 3712 2003 3715
rect 2017 3713 2019 3715
rect 2033 3713 2035 3715
rect 2038 3710 2040 3715
rect 2059 3710 2061 3715
rect 2075 3713 2077 3715
rect 2091 3713 2093 3715
rect 2096 3710 2098 3715
rect 2112 3713 2114 3715
rect 2128 3713 2130 3715
rect 2133 3712 2135 3715
rect 2149 3713 2151 3715
rect 2165 3713 2167 3715
rect 2170 3710 2172 3715
rect 2191 3710 2193 3715
rect 2207 3713 2209 3715
rect 2223 3713 2225 3715
rect 2228 3710 2230 3715
rect 2244 3713 2246 3715
rect 2260 3713 2262 3715
rect 2265 3712 2267 3715
rect 2281 3713 2283 3715
rect 2297 3713 2299 3715
rect 2302 3710 2304 3715
rect 2323 3710 2325 3715
rect 2339 3713 2341 3715
rect 2355 3713 2357 3715
rect 2360 3710 2362 3715
rect 2376 3713 2378 3715
rect 2392 3713 2394 3715
rect 2397 3712 2399 3715
rect 2413 3713 2415 3715
rect 2429 3713 2431 3715
rect 2434 3710 2436 3715
rect 2455 3710 2457 3715
rect 2471 3713 2473 3715
rect 2487 3713 2489 3715
rect 2492 3710 2494 3715
rect 2508 3713 2510 3715
rect 2589 3713 2591 3715
rect 2594 3713 2596 3716
rect 2610 3713 2612 3715
rect 2626 3713 2628 3715
rect 2631 3713 2633 3716
rect 2652 3713 2654 3716
rect 2668 3713 2670 3716
rect 2684 3713 2686 3715
rect 2689 3713 2691 3716
rect 2705 3713 2707 3715
rect 2941 3713 2943 3715
rect 2946 3712 2948 3715
rect 2962 3713 2964 3715
rect 2978 3713 2980 3715
rect 2983 3710 2985 3715
rect 3004 3710 3006 3715
rect 3020 3713 3022 3715
rect 3036 3713 3038 3715
rect 3041 3710 3043 3715
rect 3057 3713 3059 3715
rect 3073 3713 3075 3715
rect 3078 3712 3080 3715
rect 3094 3713 3096 3715
rect 3110 3713 3112 3715
rect 3115 3710 3117 3715
rect 3136 3710 3138 3715
rect 3152 3713 3154 3715
rect 3168 3713 3170 3715
rect 3173 3710 3175 3715
rect 3189 3713 3191 3715
rect 3205 3713 3207 3715
rect 3210 3712 3212 3715
rect 3226 3713 3228 3715
rect 3242 3713 3244 3715
rect 3247 3710 3249 3715
rect 3268 3710 3270 3715
rect 3284 3713 3286 3715
rect 3300 3713 3302 3715
rect 3305 3710 3307 3715
rect 3321 3713 3323 3715
rect 3337 3713 3339 3715
rect 3342 3712 3344 3715
rect 3358 3713 3360 3715
rect 3374 3713 3376 3715
rect 3379 3710 3381 3715
rect 3400 3710 3402 3715
rect 3416 3713 3418 3715
rect 3432 3713 3434 3715
rect 3437 3710 3439 3715
rect 3453 3713 3455 3715
rect 1644 3700 1646 3705
rect 1649 3703 1651 3705
rect 1644 3686 1646 3696
rect 1649 3686 1651 3693
rect 1665 3686 1667 3705
rect 1681 3696 1683 3705
rect 1686 3703 1688 3705
rect 1707 3703 1709 3705
rect 1723 3702 1725 3705
rect 1681 3686 1683 3689
rect 1686 3686 1688 3688
rect 1707 3686 1709 3688
rect 1723 3686 1725 3698
rect 1739 3696 1741 3705
rect 1744 3703 1746 3705
rect 1739 3686 1741 3689
rect 1744 3686 1746 3688
rect 1760 3686 1762 3705
rect 2589 3700 2591 3705
rect 2594 3703 2596 3705
rect 2589 3686 2591 3696
rect 2594 3686 2596 3693
rect 2610 3686 2612 3705
rect 2626 3696 2628 3705
rect 2631 3703 2633 3705
rect 2652 3703 2654 3705
rect 2668 3702 2670 3705
rect 2626 3686 2628 3689
rect 2631 3686 2633 3688
rect 2652 3686 2654 3688
rect 2668 3686 2670 3698
rect 2684 3696 2686 3705
rect 2689 3703 2691 3705
rect 2684 3686 2686 3689
rect 2689 3686 2691 3688
rect 2705 3686 2707 3705
rect 1644 3680 1646 3682
rect 1649 3679 1651 3682
rect 1665 3680 1667 3682
rect 1681 3680 1683 3682
rect 1686 3677 1688 3682
rect 1707 3677 1709 3682
rect 1723 3680 1725 3682
rect 1739 3680 1741 3682
rect 1744 3677 1746 3682
rect 1760 3680 1762 3682
rect 2589 3680 2591 3682
rect 2594 3679 2596 3682
rect 2610 3680 2612 3682
rect 2626 3680 2628 3682
rect 2175 3675 2177 3677
rect 2017 3669 2019 3672
rect 2061 3669 2063 3672
rect 2087 3669 2089 3672
rect 2133 3669 2135 3672
rect 2087 3665 2088 3669
rect 2201 3669 2203 3673
rect 2229 3675 2231 3677
rect 2256 3675 2258 3677
rect 2206 3669 2208 3672
rect 2001 3662 2003 3664
rect 2017 3662 2019 3665
rect 2033 3662 2035 3664
rect 2056 3662 2058 3664
rect 2061 3662 2063 3665
rect 2087 3662 2089 3665
rect 2108 3662 2110 3665
rect 2128 3662 2130 3664
rect 2133 3662 2135 3665
rect 2151 3662 2153 3664
rect 1768 3649 1770 3652
rect 1768 3643 1770 3645
rect 1651 3640 1653 3643
rect 2001 3640 2003 3654
rect 2017 3652 2019 3654
rect 2017 3640 2019 3642
rect 2033 3640 2035 3654
rect 2056 3649 2058 3654
rect 2061 3652 2063 3654
rect 2087 3652 2089 3654
rect 2052 3645 2058 3649
rect 2056 3640 2058 3645
rect 2061 3640 2063 3642
rect 2087 3640 2089 3642
rect 2108 3640 2110 3654
rect 2128 3649 2130 3654
rect 2133 3652 2135 3654
rect 2124 3645 2130 3649
rect 2128 3640 2130 3645
rect 2133 3640 2135 3642
rect 2151 3640 2153 3654
rect 2175 3653 2177 3667
rect 2282 3669 2284 3673
rect 2310 3675 2312 3677
rect 2631 3677 2633 3682
rect 2652 3677 2654 3682
rect 2668 3680 2670 3682
rect 2684 3680 2686 3682
rect 2689 3677 2691 3682
rect 2705 3680 2707 3682
rect 2287 3669 2289 3672
rect 2201 3658 2203 3661
rect 2206 3659 2208 3661
rect 2202 3654 2203 3658
rect 2201 3649 2203 3654
rect 2206 3649 2208 3651
rect 2175 3647 2177 3649
rect 2229 3645 2231 3667
rect 2256 3653 2258 3667
rect 3120 3675 3122 3677
rect 2282 3658 2284 3661
rect 2287 3659 2289 3661
rect 2283 3654 2284 3658
rect 2282 3649 2284 3654
rect 2287 3649 2289 3651
rect 2256 3647 2258 3649
rect 2310 3645 2312 3667
rect 2962 3669 2964 3672
rect 3006 3669 3008 3672
rect 3032 3669 3034 3672
rect 3078 3669 3080 3672
rect 3032 3665 3033 3669
rect 3146 3669 3148 3673
rect 3174 3675 3176 3677
rect 3201 3675 3203 3677
rect 3151 3669 3153 3672
rect 2946 3662 2948 3664
rect 2962 3662 2964 3665
rect 2978 3662 2980 3664
rect 3001 3662 3003 3664
rect 3006 3662 3008 3665
rect 3032 3662 3034 3665
rect 3053 3662 3055 3665
rect 3073 3662 3075 3664
rect 3078 3662 3080 3665
rect 3096 3662 3098 3664
rect 2713 3649 2715 3652
rect 2201 3643 2203 3645
rect 2206 3640 2208 3645
rect 2282 3643 2284 3645
rect 2229 3639 2231 3641
rect 2287 3640 2289 3645
rect 2713 3643 2715 3645
rect 2310 3639 2312 3641
rect 2596 3640 2598 3643
rect 2946 3640 2948 3654
rect 2962 3652 2964 3654
rect 2962 3640 2964 3642
rect 2978 3640 2980 3654
rect 3001 3649 3003 3654
rect 3006 3652 3008 3654
rect 3032 3652 3034 3654
rect 2997 3645 3003 3649
rect 3001 3640 3003 3645
rect 3006 3640 3008 3642
rect 3032 3640 3034 3642
rect 3053 3640 3055 3654
rect 3073 3649 3075 3654
rect 3078 3652 3080 3654
rect 3069 3645 3075 3649
rect 3073 3640 3075 3645
rect 3078 3640 3080 3642
rect 3096 3640 3098 3654
rect 3120 3653 3122 3667
rect 3227 3669 3229 3673
rect 3255 3675 3257 3677
rect 3232 3669 3234 3672
rect 3146 3658 3148 3661
rect 3151 3659 3153 3661
rect 3147 3654 3148 3658
rect 3146 3649 3148 3654
rect 3151 3649 3153 3651
rect 3120 3647 3122 3649
rect 3174 3645 3176 3667
rect 3201 3653 3203 3667
rect 3227 3658 3229 3661
rect 3232 3659 3234 3661
rect 3228 3654 3229 3658
rect 3227 3649 3229 3654
rect 3232 3649 3234 3651
rect 3201 3647 3203 3649
rect 3255 3645 3257 3667
rect 3146 3643 3148 3645
rect 3151 3640 3153 3645
rect 3227 3643 3229 3645
rect 3174 3639 3176 3641
rect 3232 3640 3234 3645
rect 3255 3639 3257 3641
rect 1651 3634 1653 3636
rect 2001 3634 2003 3636
rect 2017 3632 2019 3636
rect 2033 3634 2035 3636
rect 2056 3634 2058 3636
rect 2018 3628 2019 3632
rect 2061 3631 2063 3636
rect 2087 3632 2089 3636
rect 2108 3634 2110 3636
rect 2128 3634 2130 3636
rect 2017 3625 2019 3628
rect 2062 3627 2063 3631
rect 2088 3628 2089 3632
rect 2133 3631 2135 3636
rect 2151 3634 2153 3636
rect 2596 3634 2598 3636
rect 2946 3634 2948 3636
rect 2962 3632 2964 3636
rect 2978 3634 2980 3636
rect 3001 3634 3003 3636
rect 2061 3625 2063 3627
rect 2087 3624 2089 3628
rect 2134 3627 2135 3631
rect 2963 3628 2964 3632
rect 3006 3631 3008 3636
rect 3032 3632 3034 3636
rect 3053 3634 3055 3636
rect 3073 3634 3075 3636
rect 2133 3625 2135 3627
rect 2962 3625 2964 3628
rect 3007 3627 3008 3631
rect 3033 3628 3034 3632
rect 3078 3631 3080 3636
rect 3096 3634 3098 3636
rect 3006 3625 3008 3627
rect 3032 3624 3034 3628
rect 3079 3627 3080 3631
rect 3078 3625 3080 3627
rect 1635 3611 1637 3613
rect 1651 3611 1653 3614
rect 1656 3611 1658 3613
rect 1672 3611 1674 3614
rect 1688 3611 1690 3614
rect 1709 3611 1711 3614
rect 1714 3611 1716 3613
rect 1730 3611 1732 3613
rect 1746 3611 1748 3614
rect 1751 3611 1753 3613
rect 2580 3611 2582 3613
rect 2596 3611 2598 3614
rect 2601 3611 2603 3613
rect 2617 3611 2619 3614
rect 2633 3611 2635 3614
rect 2654 3611 2656 3614
rect 2659 3611 2661 3613
rect 2675 3611 2677 3613
rect 2691 3611 2693 3614
rect 2696 3611 2698 3613
rect 1635 3584 1637 3603
rect 1651 3601 1653 3603
rect 1656 3594 1658 3603
rect 1672 3600 1674 3603
rect 1688 3601 1690 3603
rect 1709 3601 1711 3603
rect 1651 3584 1653 3586
rect 1656 3584 1658 3587
rect 1672 3584 1674 3596
rect 1714 3594 1716 3603
rect 1688 3584 1690 3586
rect 1709 3584 1711 3586
rect 1714 3584 1716 3587
rect 1730 3584 1732 3603
rect 1746 3601 1748 3603
rect 1751 3598 1753 3603
rect 2017 3602 2019 3605
rect 2061 3603 2063 3605
rect 2018 3598 2019 3602
rect 2062 3599 2063 3603
rect 2087 3602 2089 3606
rect 2133 3603 2135 3605
rect 2001 3594 2003 3596
rect 2017 3594 2019 3598
rect 2033 3594 2035 3596
rect 2056 3594 2058 3596
rect 2061 3594 2063 3599
rect 2088 3598 2089 3602
rect 2134 3599 2135 3603
rect 2087 3594 2089 3598
rect 2108 3594 2110 3596
rect 2128 3594 2130 3596
rect 2133 3594 2135 3599
rect 2151 3594 2153 3596
rect 1746 3584 1748 3591
rect 1751 3584 1753 3594
rect 2201 3593 2203 3596
rect 2206 3593 2208 3596
rect 2282 3593 2284 3596
rect 2287 3593 2289 3596
rect 1635 3578 1637 3580
rect 1651 3575 1653 3580
rect 1656 3578 1658 3580
rect 1672 3578 1674 3580
rect 1688 3575 1690 3580
rect 1709 3575 1711 3580
rect 1714 3578 1716 3580
rect 1730 3578 1732 3580
rect 1746 3577 1748 3580
rect 1751 3578 1753 3580
rect 2001 3576 2003 3590
rect 2017 3588 2019 3590
rect 2017 3576 2019 3578
rect 2033 3576 2035 3590
rect 2056 3585 2058 3590
rect 2061 3588 2063 3590
rect 2087 3588 2089 3590
rect 2052 3581 2058 3585
rect 2056 3576 2058 3581
rect 2061 3576 2063 3578
rect 2087 3576 2089 3578
rect 2108 3576 2110 3590
rect 2128 3585 2130 3590
rect 2133 3588 2135 3590
rect 2124 3581 2130 3585
rect 2128 3576 2130 3581
rect 2133 3576 2135 3578
rect 2151 3576 2153 3590
rect 2201 3577 2203 3589
rect 2206 3587 2208 3589
rect 2206 3577 2208 3579
rect 2282 3577 2284 3589
rect 2287 3587 2289 3589
rect 2580 3584 2582 3603
rect 2596 3601 2598 3603
rect 2601 3594 2603 3603
rect 2617 3600 2619 3603
rect 2633 3601 2635 3603
rect 2654 3601 2656 3603
rect 2596 3584 2598 3586
rect 2601 3584 2603 3587
rect 2617 3584 2619 3596
rect 2659 3594 2661 3603
rect 2633 3584 2635 3586
rect 2654 3584 2656 3586
rect 2659 3584 2661 3587
rect 2675 3584 2677 3603
rect 2691 3601 2693 3603
rect 2696 3598 2698 3603
rect 2962 3602 2964 3605
rect 3006 3603 3008 3605
rect 2963 3598 2964 3602
rect 3007 3599 3008 3603
rect 3032 3602 3034 3606
rect 3078 3603 3080 3605
rect 2946 3594 2948 3596
rect 2962 3594 2964 3598
rect 2978 3594 2980 3596
rect 3001 3594 3003 3596
rect 3006 3594 3008 3599
rect 3033 3598 3034 3602
rect 3079 3599 3080 3603
rect 3032 3594 3034 3598
rect 3053 3594 3055 3596
rect 3073 3594 3075 3596
rect 3078 3594 3080 3599
rect 3096 3594 3098 3596
rect 2691 3584 2693 3591
rect 2696 3584 2698 3594
rect 3146 3593 3148 3596
rect 3151 3593 3153 3596
rect 3227 3593 3229 3596
rect 3232 3593 3234 3596
rect 2287 3577 2289 3579
rect 2580 3578 2582 3580
rect 2596 3575 2598 3580
rect 2601 3578 2603 3580
rect 2617 3578 2619 3580
rect 2633 3575 2635 3580
rect 2654 3575 2656 3580
rect 2659 3578 2661 3580
rect 2675 3578 2677 3580
rect 2691 3577 2693 3580
rect 2696 3578 2698 3580
rect 2946 3576 2948 3590
rect 2962 3588 2964 3590
rect 2962 3576 2964 3578
rect 2978 3576 2980 3590
rect 3001 3585 3003 3590
rect 3006 3588 3008 3590
rect 3032 3588 3034 3590
rect 2997 3581 3003 3585
rect 3001 3576 3003 3581
rect 3006 3576 3008 3578
rect 3032 3576 3034 3578
rect 3053 3576 3055 3590
rect 3073 3585 3075 3590
rect 3078 3588 3080 3590
rect 3069 3581 3075 3585
rect 3073 3576 3075 3581
rect 3078 3576 3080 3578
rect 3096 3576 3098 3590
rect 3146 3577 3148 3589
rect 3151 3587 3153 3589
rect 3151 3577 3153 3579
rect 3227 3577 3229 3589
rect 3232 3587 3234 3589
rect 3232 3577 3234 3579
rect 2001 3566 2003 3568
rect 2017 3565 2019 3568
rect 2033 3566 2035 3568
rect 2056 3566 2058 3568
rect 2061 3565 2063 3568
rect 2087 3565 2089 3568
rect 2108 3565 2110 3568
rect 2128 3566 2130 3568
rect 2133 3565 2135 3568
rect 2151 3566 2153 3568
rect 2201 3567 2203 3569
rect 2087 3561 2088 3565
rect 2206 3564 2208 3569
rect 2282 3567 2284 3569
rect 2287 3564 2289 3569
rect 2946 3566 2948 3568
rect 2962 3565 2964 3568
rect 2978 3566 2980 3568
rect 3001 3566 3003 3568
rect 3006 3565 3008 3568
rect 3032 3565 3034 3568
rect 3053 3565 3055 3568
rect 3073 3566 3075 3568
rect 3078 3565 3080 3568
rect 3096 3566 3098 3568
rect 3146 3567 3148 3569
rect 2017 3558 2019 3561
rect 2061 3558 2063 3561
rect 2087 3558 2089 3561
rect 2133 3558 2135 3561
rect 3032 3561 3033 3565
rect 3151 3564 3153 3569
rect 3227 3567 3229 3569
rect 3232 3564 3234 3569
rect 2962 3558 2964 3561
rect 3006 3558 3008 3561
rect 3032 3558 3034 3561
rect 3078 3558 3080 3561
rect 2017 3537 2019 3540
rect 2061 3537 2063 3540
rect 2087 3537 2089 3540
rect 2133 3537 2135 3540
rect 2201 3537 2203 3541
rect 2229 3543 2231 3545
rect 2280 3543 2282 3545
rect 2206 3537 2208 3540
rect 2087 3533 2088 3537
rect 2001 3530 2003 3532
rect 2017 3530 2019 3533
rect 2033 3530 2035 3532
rect 2056 3530 2058 3532
rect 2061 3530 2063 3533
rect 2087 3530 2089 3533
rect 2108 3530 2110 3533
rect 2128 3530 2130 3532
rect 2133 3530 2135 3533
rect 2151 3530 2153 3532
rect 2306 3537 2308 3541
rect 2334 3543 2336 3545
rect 2311 3537 2313 3540
rect 2201 3526 2203 3529
rect 2206 3527 2208 3529
rect 2202 3522 2203 3526
rect 2001 3508 2003 3522
rect 2017 3520 2019 3522
rect 2017 3508 2019 3510
rect 2033 3508 2035 3522
rect 2056 3517 2058 3522
rect 2061 3520 2063 3522
rect 2087 3520 2089 3522
rect 2052 3513 2058 3517
rect 2056 3508 2058 3513
rect 2061 3508 2063 3510
rect 2087 3508 2089 3510
rect 2108 3508 2110 3522
rect 2128 3517 2130 3522
rect 2133 3520 2135 3522
rect 2124 3513 2130 3517
rect 2128 3508 2130 3513
rect 2133 3508 2135 3510
rect 2151 3508 2153 3522
rect 2201 3517 2203 3522
rect 2206 3517 2208 3519
rect 2229 3513 2231 3535
rect 2280 3521 2282 3535
rect 2962 3537 2964 3540
rect 3006 3537 3008 3540
rect 3032 3537 3034 3540
rect 3078 3537 3080 3540
rect 3146 3537 3148 3541
rect 3174 3543 3176 3545
rect 3225 3543 3227 3545
rect 3151 3537 3153 3540
rect 2306 3526 2308 3529
rect 2311 3527 2313 3529
rect 2307 3522 2308 3526
rect 2306 3517 2308 3522
rect 2311 3517 2313 3519
rect 2280 3515 2282 3517
rect 2334 3513 2336 3535
rect 3032 3533 3033 3537
rect 2946 3530 2948 3532
rect 2962 3530 2964 3533
rect 2978 3530 2980 3532
rect 3001 3530 3003 3532
rect 3006 3530 3008 3533
rect 3032 3530 3034 3533
rect 3053 3530 3055 3533
rect 3073 3530 3075 3532
rect 3078 3530 3080 3533
rect 3096 3530 3098 3532
rect 3251 3537 3253 3541
rect 3279 3543 3281 3545
rect 3256 3537 3258 3540
rect 3146 3526 3148 3529
rect 3151 3527 3153 3529
rect 3147 3522 3148 3526
rect 2201 3511 2203 3513
rect 2206 3508 2208 3513
rect 2306 3511 2308 3513
rect 2229 3507 2231 3509
rect 2311 3508 2313 3513
rect 2334 3507 2336 3509
rect 2946 3508 2948 3522
rect 2962 3520 2964 3522
rect 2962 3508 2964 3510
rect 2978 3508 2980 3522
rect 3001 3517 3003 3522
rect 3006 3520 3008 3522
rect 3032 3520 3034 3522
rect 2997 3513 3003 3517
rect 3001 3508 3003 3513
rect 3006 3508 3008 3510
rect 3032 3508 3034 3510
rect 3053 3508 3055 3522
rect 3073 3517 3075 3522
rect 3078 3520 3080 3522
rect 3069 3513 3075 3517
rect 3073 3508 3075 3513
rect 3078 3508 3080 3510
rect 3096 3508 3098 3522
rect 3146 3517 3148 3522
rect 3151 3517 3153 3519
rect 3174 3513 3176 3535
rect 3225 3521 3227 3535
rect 3251 3526 3253 3529
rect 3256 3527 3258 3529
rect 3252 3522 3253 3526
rect 3251 3517 3253 3522
rect 3256 3517 3258 3519
rect 3225 3515 3227 3517
rect 3279 3513 3281 3535
rect 3146 3511 3148 3513
rect 3151 3508 3153 3513
rect 3251 3511 3253 3513
rect 3174 3507 3176 3509
rect 3256 3508 3258 3513
rect 3279 3507 3281 3509
rect 2001 3502 2003 3504
rect 2017 3500 2019 3504
rect 2033 3502 2035 3504
rect 2056 3502 2058 3504
rect 2018 3496 2019 3500
rect 2061 3499 2063 3504
rect 2087 3500 2089 3504
rect 2108 3502 2110 3504
rect 2128 3502 2130 3504
rect 2017 3493 2019 3496
rect 2062 3495 2063 3499
rect 2088 3496 2089 3500
rect 2133 3499 2135 3504
rect 2151 3502 2153 3504
rect 2946 3502 2948 3504
rect 2962 3500 2964 3504
rect 2978 3502 2980 3504
rect 3001 3502 3003 3504
rect 2061 3493 2063 3495
rect 2087 3492 2089 3496
rect 2134 3495 2135 3499
rect 2963 3496 2964 3500
rect 3006 3499 3008 3504
rect 3032 3500 3034 3504
rect 3053 3502 3055 3504
rect 3073 3502 3075 3504
rect 2133 3493 2135 3495
rect 2962 3493 2964 3496
rect 3007 3495 3008 3499
rect 3033 3496 3034 3500
rect 3078 3499 3080 3504
rect 3096 3502 3098 3504
rect 3006 3493 3008 3495
rect 3032 3492 3034 3496
rect 3079 3495 3080 3499
rect 3078 3493 3080 3495
rect 2017 3470 2019 3473
rect 2061 3471 2063 3473
rect 2018 3466 2019 3470
rect 2062 3467 2063 3471
rect 2087 3470 2089 3474
rect 2133 3471 2135 3473
rect 2001 3462 2003 3464
rect 2017 3462 2019 3466
rect 2033 3462 2035 3464
rect 2056 3462 2058 3464
rect 2061 3462 2063 3467
rect 2088 3466 2089 3470
rect 2134 3467 2135 3471
rect 2962 3470 2964 3473
rect 3006 3471 3008 3473
rect 2087 3462 2089 3466
rect 2108 3462 2110 3464
rect 2128 3462 2130 3464
rect 2133 3462 2135 3467
rect 2963 3466 2964 3470
rect 3007 3467 3008 3471
rect 3032 3470 3034 3474
rect 3078 3471 3080 3473
rect 2151 3462 2153 3464
rect 2201 3462 2203 3465
rect 2206 3462 2208 3465
rect 2306 3462 2308 3465
rect 2311 3462 2313 3465
rect 2946 3462 2948 3464
rect 2962 3462 2964 3466
rect 2978 3462 2980 3464
rect 3001 3462 3003 3464
rect 3006 3462 3008 3467
rect 3033 3466 3034 3470
rect 3079 3467 3080 3471
rect 3032 3462 3034 3466
rect 3053 3462 3055 3464
rect 3073 3462 3075 3464
rect 3078 3462 3080 3467
rect 3096 3462 3098 3464
rect 3146 3462 3148 3465
rect 3151 3462 3153 3465
rect 3251 3462 3253 3465
rect 3256 3462 3258 3465
rect 2001 3444 2003 3458
rect 2017 3456 2019 3458
rect 2017 3444 2019 3446
rect 2033 3444 2035 3458
rect 2056 3453 2058 3458
rect 2061 3456 2063 3458
rect 2087 3456 2089 3458
rect 2052 3449 2058 3453
rect 2056 3444 2058 3449
rect 2061 3444 2063 3446
rect 2087 3444 2089 3446
rect 2108 3444 2110 3458
rect 2128 3453 2130 3458
rect 2133 3456 2135 3458
rect 2124 3449 2130 3453
rect 2128 3444 2130 3449
rect 2133 3444 2135 3446
rect 2151 3444 2153 3458
rect 2201 3446 2203 3458
rect 2206 3456 2208 3458
rect 2206 3446 2208 3448
rect 2306 3446 2308 3458
rect 2311 3456 2313 3458
rect 2311 3446 2313 3448
rect 2946 3444 2948 3458
rect 2962 3456 2964 3458
rect 2962 3444 2964 3446
rect 2978 3444 2980 3458
rect 3001 3453 3003 3458
rect 3006 3456 3008 3458
rect 3032 3456 3034 3458
rect 2997 3449 3003 3453
rect 3001 3444 3003 3449
rect 3006 3444 3008 3446
rect 3032 3444 3034 3446
rect 3053 3444 3055 3458
rect 3073 3453 3075 3458
rect 3078 3456 3080 3458
rect 3069 3449 3075 3453
rect 3073 3444 3075 3449
rect 3078 3444 3080 3446
rect 3096 3444 3098 3458
rect 3146 3446 3148 3458
rect 3151 3456 3153 3458
rect 3151 3446 3153 3448
rect 3251 3446 3253 3458
rect 3256 3456 3258 3458
rect 3256 3446 3258 3448
rect 2201 3436 2203 3438
rect 2001 3434 2003 3436
rect 2017 3433 2019 3436
rect 2033 3434 2035 3436
rect 2056 3434 2058 3436
rect 2061 3433 2063 3436
rect 2087 3433 2089 3436
rect 2108 3433 2110 3436
rect 2128 3434 2130 3436
rect 2133 3433 2135 3436
rect 2151 3434 2153 3436
rect 2206 3433 2208 3438
rect 2306 3436 2308 3438
rect 2311 3433 2313 3438
rect 3146 3436 3148 3438
rect 2946 3434 2948 3436
rect 2087 3429 2088 3433
rect 2962 3433 2964 3436
rect 2978 3434 2980 3436
rect 3001 3434 3003 3436
rect 3006 3433 3008 3436
rect 3032 3433 3034 3436
rect 3053 3433 3055 3436
rect 3073 3434 3075 3436
rect 3078 3433 3080 3436
rect 3096 3434 3098 3436
rect 3151 3433 3153 3438
rect 3251 3436 3253 3438
rect 3256 3433 3258 3438
rect 3032 3429 3033 3433
rect 2017 3426 2019 3429
rect 2061 3426 2063 3429
rect 2087 3426 2089 3429
rect 2133 3426 2135 3429
rect 2962 3426 2964 3429
rect 3006 3426 3008 3429
rect 3032 3426 3034 3429
rect 3078 3426 3080 3429
rect 2017 3405 2019 3408
rect 2061 3405 2063 3408
rect 2087 3405 2089 3408
rect 2133 3405 2135 3408
rect 2201 3405 2203 3409
rect 2229 3411 2231 3413
rect 2256 3411 2258 3413
rect 2206 3405 2208 3408
rect 2087 3401 2088 3405
rect 2001 3398 2003 3400
rect 2017 3398 2019 3401
rect 2033 3398 2035 3400
rect 2056 3398 2058 3400
rect 2061 3398 2063 3401
rect 2087 3398 2089 3401
rect 2108 3398 2110 3401
rect 2128 3398 2130 3400
rect 2133 3398 2135 3401
rect 2151 3398 2153 3400
rect 2282 3405 2284 3409
rect 2310 3411 2312 3413
rect 2346 3411 2348 3413
rect 2287 3405 2289 3408
rect 2201 3394 2203 3397
rect 2206 3395 2208 3397
rect 2202 3390 2203 3394
rect 2001 3376 2003 3390
rect 2017 3388 2019 3390
rect 2017 3376 2019 3378
rect 2033 3376 2035 3390
rect 2056 3385 2058 3390
rect 2061 3388 2063 3390
rect 2087 3388 2089 3390
rect 2052 3381 2058 3385
rect 2056 3376 2058 3381
rect 2061 3376 2063 3378
rect 2087 3376 2089 3378
rect 2108 3376 2110 3390
rect 2128 3385 2130 3390
rect 2133 3388 2135 3390
rect 2124 3381 2130 3385
rect 2128 3376 2130 3381
rect 2133 3376 2135 3378
rect 2151 3376 2153 3390
rect 2201 3385 2203 3390
rect 2206 3385 2208 3387
rect 2229 3381 2231 3403
rect 2256 3389 2258 3403
rect 2372 3405 2374 3409
rect 2400 3411 2402 3413
rect 2377 3405 2379 3408
rect 2282 3394 2284 3397
rect 2287 3395 2289 3397
rect 2283 3390 2284 3394
rect 2282 3385 2284 3390
rect 2287 3385 2289 3387
rect 2256 3383 2258 3385
rect 2310 3381 2312 3403
rect 2346 3389 2348 3403
rect 2962 3405 2964 3408
rect 3006 3405 3008 3408
rect 3032 3405 3034 3408
rect 3078 3405 3080 3408
rect 3146 3405 3148 3409
rect 3174 3411 3176 3413
rect 3201 3411 3203 3413
rect 3151 3405 3153 3408
rect 2372 3394 2374 3397
rect 2377 3395 2379 3397
rect 2373 3390 2374 3394
rect 2372 3385 2374 3390
rect 2377 3385 2379 3387
rect 2346 3383 2348 3385
rect 2400 3381 2402 3403
rect 3032 3401 3033 3405
rect 2946 3398 2948 3400
rect 2962 3398 2964 3401
rect 2978 3398 2980 3400
rect 3001 3398 3003 3400
rect 3006 3398 3008 3401
rect 3032 3398 3034 3401
rect 3053 3398 3055 3401
rect 3073 3398 3075 3400
rect 3078 3398 3080 3401
rect 3096 3398 3098 3400
rect 3227 3405 3229 3409
rect 3255 3411 3257 3413
rect 3291 3411 3293 3413
rect 3232 3405 3234 3408
rect 3146 3394 3148 3397
rect 3151 3395 3153 3397
rect 3147 3390 3148 3394
rect 2201 3379 2203 3381
rect 2206 3376 2208 3381
rect 2282 3379 2284 3381
rect 2229 3375 2231 3377
rect 2287 3376 2289 3381
rect 2372 3379 2374 3381
rect 2310 3375 2312 3377
rect 2377 3376 2379 3381
rect 2400 3375 2402 3377
rect 2946 3376 2948 3390
rect 2962 3388 2964 3390
rect 2962 3376 2964 3378
rect 2978 3376 2980 3390
rect 3001 3385 3003 3390
rect 3006 3388 3008 3390
rect 3032 3388 3034 3390
rect 2997 3381 3003 3385
rect 3001 3376 3003 3381
rect 3006 3376 3008 3378
rect 3032 3376 3034 3378
rect 3053 3376 3055 3390
rect 3073 3385 3075 3390
rect 3078 3388 3080 3390
rect 3069 3381 3075 3385
rect 3073 3376 3075 3381
rect 3078 3376 3080 3378
rect 3096 3376 3098 3390
rect 3146 3385 3148 3390
rect 3151 3385 3153 3387
rect 3174 3381 3176 3403
rect 3201 3389 3203 3403
rect 3317 3405 3319 3409
rect 3345 3411 3347 3413
rect 3322 3405 3324 3408
rect 3227 3394 3229 3397
rect 3232 3395 3234 3397
rect 3228 3390 3229 3394
rect 3227 3385 3229 3390
rect 3232 3385 3234 3387
rect 3201 3383 3203 3385
rect 3255 3381 3257 3403
rect 3291 3389 3293 3403
rect 3317 3394 3319 3397
rect 3322 3395 3324 3397
rect 3318 3390 3319 3394
rect 3317 3385 3319 3390
rect 3322 3385 3324 3387
rect 3291 3383 3293 3385
rect 3345 3381 3347 3403
rect 3146 3379 3148 3381
rect 3151 3376 3153 3381
rect 3227 3379 3229 3381
rect 3174 3375 3176 3377
rect 3232 3376 3234 3381
rect 3317 3379 3319 3381
rect 3255 3375 3257 3377
rect 3322 3376 3324 3381
rect 3345 3375 3347 3377
rect 2001 3370 2003 3372
rect 2017 3368 2019 3372
rect 2033 3370 2035 3372
rect 2056 3370 2058 3372
rect 2018 3364 2019 3368
rect 2061 3367 2063 3372
rect 2087 3368 2089 3372
rect 2108 3370 2110 3372
rect 2128 3370 2130 3372
rect 2017 3361 2019 3364
rect 2062 3363 2063 3367
rect 2088 3364 2089 3368
rect 2133 3367 2135 3372
rect 2151 3370 2153 3372
rect 2946 3370 2948 3372
rect 2962 3368 2964 3372
rect 2978 3370 2980 3372
rect 3001 3370 3003 3372
rect 2061 3361 2063 3363
rect 2087 3360 2089 3364
rect 2134 3363 2135 3367
rect 2963 3364 2964 3368
rect 3006 3367 3008 3372
rect 3032 3368 3034 3372
rect 3053 3370 3055 3372
rect 3073 3370 3075 3372
rect 2133 3361 2135 3363
rect 2962 3361 2964 3364
rect 3007 3363 3008 3367
rect 3033 3364 3034 3368
rect 3078 3367 3080 3372
rect 3096 3370 3098 3372
rect 3006 3361 3008 3363
rect 3032 3360 3034 3364
rect 3079 3363 3080 3367
rect 3078 3361 3080 3363
rect 2017 3338 2019 3341
rect 2061 3339 2063 3341
rect 2018 3334 2019 3338
rect 2062 3335 2063 3339
rect 2087 3338 2089 3342
rect 2133 3339 2135 3341
rect 2001 3330 2003 3332
rect 2017 3330 2019 3334
rect 2033 3330 2035 3332
rect 2056 3330 2058 3332
rect 2061 3330 2063 3335
rect 2088 3334 2089 3338
rect 2134 3335 2135 3339
rect 2962 3338 2964 3341
rect 3006 3339 3008 3341
rect 2087 3330 2089 3334
rect 2108 3330 2110 3332
rect 2128 3330 2130 3332
rect 2133 3330 2135 3335
rect 2963 3334 2964 3338
rect 3007 3335 3008 3339
rect 3032 3338 3034 3342
rect 3078 3339 3080 3341
rect 2151 3330 2153 3332
rect 2946 3330 2948 3332
rect 2962 3330 2964 3334
rect 2978 3330 2980 3332
rect 3001 3330 3003 3332
rect 3006 3330 3008 3335
rect 3033 3334 3034 3338
rect 3079 3335 3080 3339
rect 3032 3330 3034 3334
rect 3053 3330 3055 3332
rect 3073 3330 3075 3332
rect 3078 3330 3080 3335
rect 3096 3330 3098 3332
rect 2201 3327 2203 3330
rect 2206 3327 2208 3330
rect 2282 3327 2284 3330
rect 2287 3327 2289 3330
rect 2372 3327 2374 3330
rect 2377 3327 2379 3330
rect 2001 3312 2003 3326
rect 2017 3324 2019 3326
rect 2017 3312 2019 3314
rect 2033 3312 2035 3326
rect 2056 3321 2058 3326
rect 2061 3324 2063 3326
rect 2087 3324 2089 3326
rect 2052 3317 2058 3321
rect 2056 3312 2058 3317
rect 2061 3312 2063 3314
rect 2087 3312 2089 3314
rect 2108 3312 2110 3326
rect 2128 3321 2130 3326
rect 2133 3324 2135 3326
rect 2124 3317 2130 3321
rect 2128 3312 2130 3317
rect 2133 3312 2135 3314
rect 2151 3312 2153 3326
rect 3146 3327 3148 3330
rect 3151 3327 3153 3330
rect 3227 3327 3229 3330
rect 3232 3327 3234 3330
rect 3317 3327 3319 3330
rect 3322 3327 3324 3330
rect 2201 3311 2203 3323
rect 2206 3321 2208 3323
rect 2206 3311 2208 3313
rect 2282 3311 2284 3323
rect 2287 3321 2289 3323
rect 2287 3311 2289 3313
rect 2372 3311 2374 3323
rect 2377 3321 2379 3323
rect 2377 3311 2379 3313
rect 2946 3312 2948 3326
rect 2962 3324 2964 3326
rect 2962 3312 2964 3314
rect 2978 3312 2980 3326
rect 3001 3321 3003 3326
rect 3006 3324 3008 3326
rect 3032 3324 3034 3326
rect 2997 3317 3003 3321
rect 3001 3312 3003 3317
rect 3006 3312 3008 3314
rect 3032 3312 3034 3314
rect 3053 3312 3055 3326
rect 3073 3321 3075 3326
rect 3078 3324 3080 3326
rect 3069 3317 3075 3321
rect 3073 3312 3075 3317
rect 3078 3312 3080 3314
rect 3096 3312 3098 3326
rect 2001 3302 2003 3304
rect 2017 3301 2019 3304
rect 2033 3302 2035 3304
rect 2056 3302 2058 3304
rect 2061 3301 2063 3304
rect 2087 3301 2089 3304
rect 2108 3301 2110 3304
rect 2128 3302 2130 3304
rect 2133 3301 2135 3304
rect 2151 3302 2153 3304
rect 3146 3311 3148 3323
rect 3151 3321 3153 3323
rect 3151 3311 3153 3313
rect 3227 3311 3229 3323
rect 3232 3321 3234 3323
rect 3232 3311 3234 3313
rect 3317 3311 3319 3323
rect 3322 3321 3324 3323
rect 3322 3311 3324 3313
rect 2201 3301 2203 3303
rect 2087 3297 2088 3301
rect 2206 3298 2208 3303
rect 2282 3301 2284 3303
rect 2287 3298 2289 3303
rect 2372 3301 2374 3303
rect 2377 3298 2379 3303
rect 2946 3302 2948 3304
rect 2017 3294 2019 3297
rect 2061 3294 2063 3297
rect 2087 3294 2089 3297
rect 2133 3294 2135 3297
rect 2962 3301 2964 3304
rect 2978 3302 2980 3304
rect 3001 3302 3003 3304
rect 3006 3301 3008 3304
rect 3032 3301 3034 3304
rect 3053 3301 3055 3304
rect 3073 3302 3075 3304
rect 3078 3301 3080 3304
rect 3096 3302 3098 3304
rect 3146 3301 3148 3303
rect 3032 3297 3033 3301
rect 3151 3298 3153 3303
rect 3227 3301 3229 3303
rect 3232 3298 3234 3303
rect 3317 3301 3319 3303
rect 3322 3298 3324 3303
rect 2962 3294 2964 3297
rect 3006 3294 3008 3297
rect 3032 3294 3034 3297
rect 3078 3294 3080 3297
rect 2017 3273 2019 3276
rect 2061 3273 2063 3276
rect 2087 3273 2089 3276
rect 2133 3273 2135 3276
rect 2201 3273 2203 3277
rect 2229 3279 2231 3281
rect 2206 3273 2208 3276
rect 2087 3269 2088 3273
rect 2001 3266 2003 3268
rect 2017 3266 2019 3269
rect 2033 3266 2035 3268
rect 2056 3266 2058 3268
rect 2061 3266 2063 3269
rect 2087 3266 2089 3269
rect 2108 3266 2110 3269
rect 2128 3266 2130 3268
rect 2133 3266 2135 3269
rect 2151 3266 2153 3268
rect 2962 3273 2964 3276
rect 3006 3273 3008 3276
rect 3032 3273 3034 3276
rect 3078 3273 3080 3276
rect 3146 3273 3148 3277
rect 3174 3279 3176 3281
rect 3151 3273 3153 3276
rect 2201 3262 2203 3265
rect 2206 3263 2208 3265
rect 2202 3258 2203 3262
rect 2001 3244 2003 3258
rect 2017 3256 2019 3258
rect 2017 3244 2019 3246
rect 2033 3244 2035 3258
rect 2056 3253 2058 3258
rect 2061 3256 2063 3258
rect 2087 3256 2089 3258
rect 2052 3249 2058 3253
rect 2056 3244 2058 3249
rect 2061 3244 2063 3246
rect 2087 3244 2089 3246
rect 2108 3244 2110 3258
rect 2128 3253 2130 3258
rect 2133 3256 2135 3258
rect 2124 3249 2130 3253
rect 2128 3244 2130 3249
rect 2133 3244 2135 3246
rect 2151 3244 2153 3258
rect 2201 3253 2203 3258
rect 2206 3253 2208 3255
rect 2229 3249 2231 3271
rect 3032 3269 3033 3273
rect 2946 3266 2948 3268
rect 2962 3266 2964 3269
rect 2978 3266 2980 3268
rect 3001 3266 3003 3268
rect 3006 3266 3008 3269
rect 3032 3266 3034 3269
rect 3053 3266 3055 3269
rect 3073 3266 3075 3268
rect 3078 3266 3080 3269
rect 3096 3266 3098 3268
rect 3146 3262 3148 3265
rect 3151 3263 3153 3265
rect 3147 3258 3148 3262
rect 2201 3247 2203 3249
rect 2206 3244 2208 3249
rect 2229 3243 2231 3245
rect 2946 3244 2948 3258
rect 2962 3256 2964 3258
rect 2962 3244 2964 3246
rect 2978 3244 2980 3258
rect 3001 3253 3003 3258
rect 3006 3256 3008 3258
rect 3032 3256 3034 3258
rect 2997 3249 3003 3253
rect 3001 3244 3003 3249
rect 3006 3244 3008 3246
rect 3032 3244 3034 3246
rect 3053 3244 3055 3258
rect 3073 3253 3075 3258
rect 3078 3256 3080 3258
rect 3069 3249 3075 3253
rect 3073 3244 3075 3249
rect 3078 3244 3080 3246
rect 3096 3244 3098 3258
rect 3146 3253 3148 3258
rect 3151 3253 3153 3255
rect 3174 3249 3176 3271
rect 3146 3247 3148 3249
rect 3151 3244 3153 3249
rect 3174 3243 3176 3245
rect 2001 3238 2003 3240
rect 2017 3236 2019 3240
rect 2033 3238 2035 3240
rect 2056 3238 2058 3240
rect 2018 3232 2019 3236
rect 2061 3235 2063 3240
rect 2087 3236 2089 3240
rect 2108 3238 2110 3240
rect 2128 3238 2130 3240
rect 2017 3229 2019 3232
rect 2062 3231 2063 3235
rect 2088 3232 2089 3236
rect 2133 3235 2135 3240
rect 2151 3238 2153 3240
rect 2946 3238 2948 3240
rect 2962 3236 2964 3240
rect 2978 3238 2980 3240
rect 3001 3238 3003 3240
rect 2061 3229 2063 3231
rect 2087 3228 2089 3232
rect 2134 3231 2135 3235
rect 2963 3232 2964 3236
rect 3006 3235 3008 3240
rect 3032 3236 3034 3240
rect 3053 3238 3055 3240
rect 3073 3238 3075 3240
rect 2133 3229 2135 3231
rect 2962 3229 2964 3232
rect 3007 3231 3008 3235
rect 3033 3232 3034 3236
rect 3078 3235 3080 3240
rect 3096 3238 3098 3240
rect 3006 3229 3008 3231
rect 3032 3228 3034 3232
rect 3079 3231 3080 3235
rect 3078 3229 3080 3231
rect 1512 3211 1514 3213
rect 1517 3211 1519 3214
rect 1533 3211 1535 3213
rect 1549 3211 1551 3213
rect 1554 3211 1556 3214
rect 1575 3211 1577 3214
rect 1591 3211 1593 3214
rect 1607 3211 1609 3213
rect 1612 3211 1614 3214
rect 1628 3211 1630 3213
rect 1644 3211 1646 3213
rect 1649 3211 1651 3214
rect 1665 3211 1667 3213
rect 1681 3211 1683 3213
rect 1686 3211 1688 3214
rect 1707 3211 1709 3214
rect 1723 3211 1725 3214
rect 1739 3211 1741 3213
rect 1744 3211 1746 3214
rect 1760 3211 1762 3213
rect 1776 3211 1778 3213
rect 1781 3211 1783 3214
rect 1797 3211 1799 3213
rect 1813 3211 1815 3213
rect 1818 3211 1820 3214
rect 1839 3211 1841 3214
rect 1855 3211 1857 3214
rect 1871 3211 1873 3213
rect 1876 3211 1878 3214
rect 1892 3211 1894 3213
rect 2457 3211 2459 3213
rect 2462 3211 2464 3214
rect 2478 3211 2480 3213
rect 2494 3211 2496 3213
rect 2499 3211 2501 3214
rect 2520 3211 2522 3214
rect 2536 3211 2538 3214
rect 2552 3211 2554 3213
rect 2557 3211 2559 3214
rect 2573 3211 2575 3213
rect 2589 3211 2591 3213
rect 2594 3211 2596 3214
rect 2610 3211 2612 3213
rect 2626 3211 2628 3213
rect 2631 3211 2633 3214
rect 2652 3211 2654 3214
rect 2668 3211 2670 3214
rect 2684 3211 2686 3213
rect 2689 3211 2691 3214
rect 2705 3211 2707 3213
rect 2721 3211 2723 3213
rect 2726 3211 2728 3214
rect 2742 3211 2744 3213
rect 2758 3211 2760 3213
rect 2763 3211 2765 3214
rect 2784 3211 2786 3214
rect 2800 3211 2802 3214
rect 2816 3211 2818 3213
rect 2821 3211 2823 3214
rect 2837 3211 2839 3213
rect 2017 3206 2019 3209
rect 2061 3207 2063 3209
rect 1512 3198 1514 3203
rect 1517 3201 1519 3203
rect 1512 3184 1514 3194
rect 1517 3184 1519 3191
rect 1533 3184 1535 3203
rect 1549 3194 1551 3203
rect 1554 3201 1556 3203
rect 1575 3201 1577 3203
rect 1591 3200 1593 3203
rect 1549 3184 1551 3187
rect 1554 3184 1556 3186
rect 1575 3184 1577 3186
rect 1591 3184 1593 3196
rect 1607 3194 1609 3203
rect 1612 3201 1614 3203
rect 1607 3184 1609 3187
rect 1612 3184 1614 3186
rect 1628 3184 1630 3203
rect 1644 3200 1646 3203
rect 1649 3201 1651 3203
rect 1644 3184 1646 3196
rect 1649 3184 1651 3191
rect 1665 3184 1667 3203
rect 1681 3194 1683 3203
rect 1686 3201 1688 3203
rect 1707 3201 1709 3203
rect 1723 3200 1725 3203
rect 1681 3184 1683 3187
rect 1686 3184 1688 3186
rect 1707 3184 1709 3186
rect 1723 3184 1725 3196
rect 1739 3194 1741 3203
rect 1744 3201 1746 3203
rect 1739 3184 1741 3187
rect 1744 3184 1746 3186
rect 1760 3184 1762 3203
rect 1776 3200 1778 3203
rect 1781 3201 1783 3203
rect 1776 3184 1778 3196
rect 1781 3184 1783 3191
rect 1797 3184 1799 3203
rect 1813 3194 1815 3203
rect 1818 3201 1820 3203
rect 1839 3201 1841 3203
rect 1855 3200 1857 3203
rect 1813 3184 1815 3187
rect 1818 3184 1820 3186
rect 1839 3184 1841 3186
rect 1855 3184 1857 3196
rect 1871 3194 1873 3203
rect 1876 3201 1878 3203
rect 1892 3195 1894 3203
rect 2018 3202 2019 3206
rect 2062 3203 2063 3207
rect 2087 3206 2089 3210
rect 2133 3207 2135 3209
rect 2001 3198 2003 3200
rect 2017 3198 2019 3202
rect 2033 3198 2035 3200
rect 2056 3198 2058 3200
rect 2061 3198 2063 3203
rect 2088 3202 2089 3206
rect 2134 3203 2135 3207
rect 2278 3206 2280 3209
rect 2322 3207 2324 3209
rect 2087 3198 2089 3202
rect 2108 3198 2110 3200
rect 2128 3198 2130 3200
rect 2133 3198 2135 3203
rect 2279 3202 2280 3206
rect 2323 3203 2324 3207
rect 2348 3206 2350 3210
rect 2394 3207 2396 3209
rect 2151 3198 2153 3200
rect 2235 3198 2237 3201
rect 2253 3198 2255 3201
rect 2278 3198 2280 3202
rect 2294 3198 2296 3200
rect 2317 3198 2319 3200
rect 2322 3198 2324 3203
rect 2349 3202 2350 3206
rect 2395 3203 2396 3207
rect 2962 3206 2964 3209
rect 3006 3207 3008 3209
rect 2348 3198 2350 3202
rect 2369 3198 2371 3200
rect 2389 3198 2391 3200
rect 2394 3198 2396 3203
rect 2412 3198 2414 3200
rect 2457 3198 2459 3203
rect 2462 3201 2464 3203
rect 1871 3184 1873 3187
rect 1876 3184 1878 3186
rect 1892 3184 1894 3191
rect 2001 3180 2003 3194
rect 2017 3192 2019 3194
rect 2017 3180 2019 3182
rect 2033 3180 2035 3194
rect 2056 3189 2058 3194
rect 2061 3192 2063 3194
rect 2087 3192 2089 3194
rect 2052 3185 2058 3189
rect 2056 3180 2058 3185
rect 2061 3180 2063 3182
rect 2087 3180 2089 3182
rect 2108 3180 2110 3194
rect 2128 3189 2130 3194
rect 2133 3192 2135 3194
rect 2124 3185 2130 3189
rect 2128 3180 2130 3185
rect 2133 3180 2135 3182
rect 2151 3180 2153 3194
rect 2201 3191 2203 3194
rect 2206 3191 2208 3194
rect 2235 3189 2237 3194
rect 1512 3178 1514 3180
rect 1517 3177 1519 3180
rect 1533 3178 1535 3180
rect 1549 3178 1551 3180
rect 1554 3175 1556 3180
rect 1575 3175 1577 3180
rect 1591 3178 1593 3180
rect 1607 3178 1609 3180
rect 1612 3175 1614 3180
rect 1628 3178 1630 3180
rect 1644 3178 1646 3180
rect 1649 3177 1651 3180
rect 1665 3178 1667 3180
rect 1681 3178 1683 3180
rect 1686 3175 1688 3180
rect 1707 3175 1709 3180
rect 1723 3178 1725 3180
rect 1739 3178 1741 3180
rect 1744 3175 1746 3180
rect 1760 3178 1762 3180
rect 1776 3178 1778 3180
rect 1781 3177 1783 3180
rect 1797 3178 1799 3180
rect 1813 3178 1815 3180
rect 1818 3175 1820 3180
rect 1839 3175 1841 3180
rect 1855 3178 1857 3180
rect 1871 3178 1873 3180
rect 1876 3175 1878 3180
rect 1892 3178 1894 3180
rect 2201 3175 2203 3187
rect 2206 3185 2208 3187
rect 2235 3180 2237 3185
rect 2253 3180 2255 3194
rect 2278 3192 2280 3194
rect 2278 3180 2280 3182
rect 2294 3180 2296 3194
rect 2317 3189 2319 3194
rect 2322 3192 2324 3194
rect 2348 3192 2350 3194
rect 2313 3185 2319 3189
rect 2317 3180 2319 3185
rect 2322 3180 2324 3182
rect 2348 3180 2350 3182
rect 2369 3180 2371 3194
rect 2389 3189 2391 3194
rect 2394 3192 2396 3194
rect 2385 3185 2391 3189
rect 2389 3180 2391 3185
rect 2394 3180 2396 3182
rect 2412 3180 2414 3194
rect 2457 3184 2459 3194
rect 2462 3184 2464 3191
rect 2478 3184 2480 3203
rect 2494 3194 2496 3203
rect 2499 3201 2501 3203
rect 2520 3201 2522 3203
rect 2536 3200 2538 3203
rect 2494 3184 2496 3187
rect 2499 3184 2501 3186
rect 2520 3184 2522 3186
rect 2536 3184 2538 3196
rect 2552 3194 2554 3203
rect 2557 3201 2559 3203
rect 2552 3184 2554 3187
rect 2557 3184 2559 3186
rect 2573 3184 2575 3203
rect 2589 3200 2591 3203
rect 2594 3201 2596 3203
rect 2589 3184 2591 3196
rect 2594 3184 2596 3191
rect 2610 3184 2612 3203
rect 2626 3194 2628 3203
rect 2631 3201 2633 3203
rect 2652 3201 2654 3203
rect 2668 3200 2670 3203
rect 2626 3184 2628 3187
rect 2631 3184 2633 3186
rect 2652 3184 2654 3186
rect 2668 3184 2670 3196
rect 2684 3194 2686 3203
rect 2689 3201 2691 3203
rect 2684 3184 2686 3187
rect 2689 3184 2691 3186
rect 2705 3184 2707 3203
rect 2721 3200 2723 3203
rect 2726 3201 2728 3203
rect 2721 3184 2723 3196
rect 2726 3184 2728 3191
rect 2742 3184 2744 3203
rect 2758 3194 2760 3203
rect 2763 3201 2765 3203
rect 2784 3201 2786 3203
rect 2800 3200 2802 3203
rect 2758 3184 2760 3187
rect 2763 3184 2765 3186
rect 2784 3184 2786 3186
rect 2800 3184 2802 3196
rect 2816 3194 2818 3203
rect 2821 3201 2823 3203
rect 2837 3195 2839 3203
rect 2963 3202 2964 3206
rect 3007 3203 3008 3207
rect 3032 3206 3034 3210
rect 3078 3207 3080 3209
rect 2946 3198 2948 3200
rect 2962 3198 2964 3202
rect 2978 3198 2980 3200
rect 3001 3198 3003 3200
rect 3006 3198 3008 3203
rect 3033 3202 3034 3206
rect 3079 3203 3080 3207
rect 3223 3206 3225 3209
rect 3267 3207 3269 3209
rect 3032 3198 3034 3202
rect 3053 3198 3055 3200
rect 3073 3198 3075 3200
rect 3078 3198 3080 3203
rect 3224 3202 3225 3206
rect 3268 3203 3269 3207
rect 3293 3206 3295 3210
rect 3339 3207 3341 3209
rect 3096 3198 3098 3200
rect 3180 3198 3182 3201
rect 3198 3198 3200 3201
rect 3223 3198 3225 3202
rect 3239 3198 3241 3200
rect 3262 3198 3264 3200
rect 3267 3198 3269 3203
rect 3294 3202 3295 3206
rect 3340 3203 3341 3207
rect 3293 3198 3295 3202
rect 3314 3198 3316 3200
rect 3334 3198 3336 3200
rect 3339 3198 3341 3203
rect 3357 3198 3359 3200
rect 2816 3184 2818 3187
rect 2821 3184 2823 3186
rect 2837 3184 2839 3191
rect 2946 3180 2948 3194
rect 2962 3192 2964 3194
rect 2962 3180 2964 3182
rect 2978 3180 2980 3194
rect 3001 3189 3003 3194
rect 3006 3192 3008 3194
rect 3032 3192 3034 3194
rect 2997 3185 3003 3189
rect 3001 3180 3003 3185
rect 3006 3180 3008 3182
rect 3032 3180 3034 3182
rect 3053 3180 3055 3194
rect 3073 3189 3075 3194
rect 3078 3192 3080 3194
rect 3069 3185 3075 3189
rect 3073 3180 3075 3185
rect 3078 3180 3080 3182
rect 3096 3180 3098 3194
rect 3146 3191 3148 3194
rect 3151 3191 3153 3194
rect 3180 3189 3182 3194
rect 2206 3175 2208 3177
rect 2001 3170 2003 3172
rect 2017 3169 2019 3172
rect 2033 3170 2035 3172
rect 2056 3170 2058 3172
rect 2061 3169 2063 3172
rect 2087 3169 2089 3172
rect 2108 3169 2110 3172
rect 2128 3170 2130 3172
rect 2133 3169 2135 3172
rect 2151 3170 2153 3172
rect 2087 3165 2088 3169
rect 2457 3178 2459 3180
rect 2462 3177 2464 3180
rect 2478 3178 2480 3180
rect 2494 3178 2496 3180
rect 2499 3175 2501 3180
rect 2520 3175 2522 3180
rect 2536 3178 2538 3180
rect 2552 3178 2554 3180
rect 2557 3175 2559 3180
rect 2573 3178 2575 3180
rect 2589 3178 2591 3180
rect 2235 3169 2237 3172
rect 2201 3165 2203 3167
rect 2017 3162 2019 3165
rect 2061 3162 2063 3165
rect 2087 3162 2089 3165
rect 2133 3162 2135 3165
rect 2206 3162 2208 3167
rect 1627 3140 1629 3143
rect 1651 3140 1653 3143
rect 1627 3133 1629 3136
rect 1651 3133 1653 3136
rect 2253 3130 2255 3172
rect 2278 3169 2280 3172
rect 2294 3170 2296 3172
rect 2317 3170 2319 3172
rect 2322 3169 2324 3172
rect 2348 3169 2350 3172
rect 2369 3169 2371 3172
rect 2389 3170 2391 3172
rect 2394 3169 2396 3172
rect 2412 3170 2414 3172
rect 2594 3177 2596 3180
rect 2610 3178 2612 3180
rect 2626 3178 2628 3180
rect 2631 3175 2633 3180
rect 2652 3175 2654 3180
rect 2668 3178 2670 3180
rect 2684 3178 2686 3180
rect 2689 3175 2691 3180
rect 2705 3178 2707 3180
rect 2721 3178 2723 3180
rect 2726 3177 2728 3180
rect 2742 3178 2744 3180
rect 2758 3178 2760 3180
rect 2763 3175 2765 3180
rect 2784 3175 2786 3180
rect 2800 3178 2802 3180
rect 2816 3178 2818 3180
rect 2821 3175 2823 3180
rect 2837 3178 2839 3180
rect 3146 3175 3148 3187
rect 3151 3185 3153 3187
rect 3180 3180 3182 3185
rect 3198 3180 3200 3194
rect 3223 3192 3225 3194
rect 3223 3180 3225 3182
rect 3239 3180 3241 3194
rect 3262 3189 3264 3194
rect 3267 3192 3269 3194
rect 3293 3192 3295 3194
rect 3258 3185 3264 3189
rect 3262 3180 3264 3185
rect 3267 3180 3269 3182
rect 3293 3180 3295 3182
rect 3314 3180 3316 3194
rect 3334 3189 3336 3194
rect 3339 3192 3341 3194
rect 3330 3185 3336 3189
rect 3334 3180 3336 3185
rect 3339 3180 3341 3182
rect 3357 3180 3359 3194
rect 3151 3175 3153 3177
rect 2946 3170 2948 3172
rect 2962 3169 2964 3172
rect 2978 3170 2980 3172
rect 3001 3170 3003 3172
rect 3006 3169 3008 3172
rect 3032 3169 3034 3172
rect 3053 3169 3055 3172
rect 3073 3170 3075 3172
rect 3078 3169 3080 3172
rect 3096 3170 3098 3172
rect 2348 3165 2349 3169
rect 2278 3162 2280 3165
rect 2322 3162 2324 3165
rect 2348 3162 2350 3165
rect 2394 3162 2396 3165
rect 3032 3165 3033 3169
rect 3180 3169 3182 3172
rect 3146 3165 3148 3167
rect 2962 3162 2964 3165
rect 3006 3162 3008 3165
rect 3032 3162 3034 3165
rect 3078 3162 3080 3165
rect 3151 3162 3153 3167
rect 2572 3140 2574 3143
rect 2596 3140 2598 3143
rect 2421 3138 2424 3140
rect 2428 3138 2431 3140
rect 2572 3133 2574 3136
rect 2596 3133 2598 3136
rect 3198 3134 3200 3172
rect 3223 3169 3225 3172
rect 3239 3170 3241 3172
rect 3262 3170 3264 3172
rect 3267 3169 3269 3172
rect 3293 3169 3295 3172
rect 3314 3169 3316 3172
rect 3334 3170 3336 3172
rect 3339 3169 3341 3172
rect 3357 3170 3359 3172
rect 3293 3165 3294 3169
rect 3223 3162 3225 3165
rect 3267 3162 3269 3165
rect 3293 3162 3295 3165
rect 3339 3162 3341 3165
rect 3366 3138 3369 3140
rect 3373 3138 3376 3140
rect 1647 3127 1649 3129
rect 2592 3127 2594 3129
rect 1647 3120 1649 3123
rect 2592 3120 2594 3123
rect 1636 3109 1638 3111
rect 1642 3109 1661 3111
rect 2581 3109 2583 3111
rect 2587 3109 2606 3111
rect 1627 3104 1629 3106
rect 1651 3104 1653 3106
rect 2572 3104 2574 3106
rect 2596 3104 2598 3106
rect 1627 3097 1629 3100
rect 1651 3097 1653 3100
rect 2295 3099 2297 3101
rect 2300 3099 2302 3102
rect 2316 3099 2318 3101
rect 2332 3099 2334 3101
rect 2337 3099 2339 3102
rect 2358 3099 2360 3102
rect 2374 3099 2376 3102
rect 2390 3099 2392 3101
rect 2395 3099 2397 3102
rect 2411 3099 2413 3101
rect 2572 3097 2574 3100
rect 2596 3097 2598 3100
rect 3240 3099 3242 3101
rect 3245 3099 3247 3102
rect 3261 3099 3263 3101
rect 3277 3099 3279 3101
rect 3282 3099 3284 3102
rect 3303 3099 3305 3102
rect 3319 3099 3321 3102
rect 3335 3099 3337 3101
rect 3340 3099 3342 3102
rect 3356 3099 3358 3101
rect 2295 3086 2297 3091
rect 2300 3089 2302 3091
rect 2295 3072 2297 3082
rect 2300 3072 2302 3079
rect 2316 3072 2318 3091
rect 2332 3082 2334 3091
rect 2337 3089 2339 3091
rect 2358 3089 2360 3091
rect 2374 3088 2376 3091
rect 2332 3072 2334 3075
rect 2337 3072 2339 3074
rect 2358 3072 2360 3074
rect 2374 3072 2376 3084
rect 2390 3082 2392 3091
rect 2395 3089 2397 3091
rect 2390 3072 2392 3075
rect 2395 3072 2397 3074
rect 2411 3072 2413 3091
rect 3240 3086 3242 3091
rect 3245 3089 3247 3091
rect 3240 3072 3242 3082
rect 3245 3072 3247 3079
rect 3261 3072 3263 3091
rect 3277 3082 3279 3091
rect 3282 3089 3284 3091
rect 3303 3089 3305 3091
rect 3319 3088 3321 3091
rect 3277 3072 3279 3075
rect 3282 3072 3284 3074
rect 3303 3072 3305 3074
rect 3319 3072 3321 3084
rect 3335 3082 3337 3091
rect 3340 3089 3342 3091
rect 3335 3072 3337 3075
rect 3340 3072 3342 3074
rect 3356 3072 3358 3091
rect 1512 3069 1514 3071
rect 1517 3069 1519 3072
rect 1533 3069 1535 3071
rect 1549 3069 1551 3071
rect 1554 3069 1556 3072
rect 1575 3069 1577 3072
rect 1591 3069 1593 3072
rect 1607 3069 1609 3071
rect 1612 3069 1614 3072
rect 1628 3069 1630 3071
rect 1644 3069 1646 3071
rect 1649 3069 1651 3072
rect 1665 3069 1667 3071
rect 1681 3069 1683 3071
rect 1686 3069 1688 3072
rect 1707 3069 1709 3072
rect 1723 3069 1725 3072
rect 1739 3069 1741 3071
rect 1744 3069 1746 3072
rect 1760 3069 1762 3071
rect 1776 3069 1778 3071
rect 1781 3069 1783 3072
rect 1797 3069 1799 3071
rect 1813 3069 1815 3071
rect 1818 3069 1820 3072
rect 1839 3069 1841 3072
rect 1855 3069 1857 3072
rect 1871 3069 1873 3071
rect 1876 3069 1878 3072
rect 1892 3069 1894 3071
rect 2457 3069 2459 3071
rect 2462 3069 2464 3072
rect 2478 3069 2480 3071
rect 2494 3069 2496 3071
rect 2499 3069 2501 3072
rect 2520 3069 2522 3072
rect 2536 3069 2538 3072
rect 2552 3069 2554 3071
rect 2557 3069 2559 3072
rect 2573 3069 2575 3071
rect 2589 3069 2591 3071
rect 2594 3069 2596 3072
rect 2610 3069 2612 3071
rect 2626 3069 2628 3071
rect 2631 3069 2633 3072
rect 2652 3069 2654 3072
rect 2668 3069 2670 3072
rect 2684 3069 2686 3071
rect 2689 3069 2691 3072
rect 2705 3069 2707 3071
rect 2721 3069 2723 3071
rect 2726 3069 2728 3072
rect 2742 3069 2744 3071
rect 2758 3069 2760 3071
rect 2763 3069 2765 3072
rect 2784 3069 2786 3072
rect 2800 3069 2802 3072
rect 2816 3069 2818 3071
rect 2821 3069 2823 3072
rect 2837 3069 2839 3071
rect 2295 3066 2297 3068
rect 2300 3065 2302 3068
rect 2316 3066 2318 3068
rect 2332 3066 2334 3068
rect 2337 3063 2339 3068
rect 2358 3063 2360 3068
rect 2374 3066 2376 3068
rect 2390 3066 2392 3068
rect 2395 3063 2397 3068
rect 2411 3066 2413 3068
rect 1512 3056 1514 3061
rect 1517 3059 1519 3061
rect 1512 3042 1514 3052
rect 1517 3042 1519 3049
rect 1533 3042 1535 3061
rect 1549 3052 1551 3061
rect 1554 3059 1556 3061
rect 1575 3059 1577 3061
rect 1591 3058 1593 3061
rect 1549 3042 1551 3045
rect 1554 3042 1556 3044
rect 1575 3042 1577 3044
rect 1591 3042 1593 3054
rect 1607 3052 1609 3061
rect 1612 3059 1614 3061
rect 1607 3042 1609 3045
rect 1612 3042 1614 3044
rect 1628 3042 1630 3061
rect 1644 3058 1646 3061
rect 1649 3059 1651 3061
rect 1644 3042 1646 3054
rect 1649 3042 1651 3049
rect 1665 3042 1667 3061
rect 1681 3052 1683 3061
rect 1686 3059 1688 3061
rect 1707 3059 1709 3061
rect 1723 3058 1725 3061
rect 1681 3042 1683 3045
rect 1686 3042 1688 3044
rect 1707 3042 1709 3044
rect 1723 3042 1725 3054
rect 1739 3052 1741 3061
rect 1744 3059 1746 3061
rect 1739 3042 1741 3045
rect 1744 3042 1746 3044
rect 1760 3042 1762 3061
rect 1776 3058 1778 3061
rect 1781 3059 1783 3061
rect 1776 3042 1778 3054
rect 1781 3042 1783 3049
rect 1797 3042 1799 3061
rect 1813 3052 1815 3061
rect 1818 3059 1820 3061
rect 1839 3059 1841 3061
rect 1855 3058 1857 3061
rect 1813 3042 1815 3045
rect 1818 3042 1820 3044
rect 1839 3042 1841 3044
rect 1855 3042 1857 3054
rect 1871 3052 1873 3061
rect 1876 3059 1878 3061
rect 1892 3053 1894 3061
rect 3240 3066 3242 3068
rect 3245 3065 3247 3068
rect 3261 3066 3263 3068
rect 3277 3066 3279 3068
rect 3282 3063 3284 3068
rect 3303 3063 3305 3068
rect 3319 3066 3321 3068
rect 3335 3066 3337 3068
rect 3340 3063 3342 3068
rect 3356 3066 3358 3068
rect 2457 3056 2459 3061
rect 2462 3059 2464 3061
rect 1871 3042 1873 3045
rect 1876 3042 1878 3044
rect 1892 3042 1894 3049
rect 2457 3042 2459 3052
rect 2462 3042 2464 3049
rect 2478 3042 2480 3061
rect 2494 3052 2496 3061
rect 2499 3059 2501 3061
rect 2520 3059 2522 3061
rect 2536 3058 2538 3061
rect 2494 3042 2496 3045
rect 2499 3042 2501 3044
rect 2520 3042 2522 3044
rect 2536 3042 2538 3054
rect 2552 3052 2554 3061
rect 2557 3059 2559 3061
rect 2552 3042 2554 3045
rect 2557 3042 2559 3044
rect 2573 3042 2575 3061
rect 2589 3058 2591 3061
rect 2594 3059 2596 3061
rect 2589 3042 2591 3054
rect 2594 3042 2596 3049
rect 2610 3042 2612 3061
rect 2626 3052 2628 3061
rect 2631 3059 2633 3061
rect 2652 3059 2654 3061
rect 2668 3058 2670 3061
rect 2626 3042 2628 3045
rect 2631 3042 2633 3044
rect 2652 3042 2654 3044
rect 2668 3042 2670 3054
rect 2684 3052 2686 3061
rect 2689 3059 2691 3061
rect 2684 3042 2686 3045
rect 2689 3042 2691 3044
rect 2705 3042 2707 3061
rect 2721 3058 2723 3061
rect 2726 3059 2728 3061
rect 2721 3042 2723 3054
rect 2726 3042 2728 3049
rect 2742 3042 2744 3061
rect 2758 3052 2760 3061
rect 2763 3059 2765 3061
rect 2784 3059 2786 3061
rect 2800 3058 2802 3061
rect 2758 3042 2760 3045
rect 2763 3042 2765 3044
rect 2784 3042 2786 3044
rect 2800 3042 2802 3054
rect 2816 3052 2818 3061
rect 2821 3059 2823 3061
rect 2837 3053 2839 3061
rect 2816 3042 2818 3045
rect 2821 3042 2823 3044
rect 2837 3042 2839 3049
rect 1512 3036 1514 3038
rect 1517 3035 1519 3038
rect 1533 3036 1535 3038
rect 1549 3036 1551 3038
rect 1554 3033 1556 3038
rect 1575 3033 1577 3038
rect 1591 3036 1593 3038
rect 1607 3036 1609 3038
rect 1612 3033 1614 3038
rect 1628 3036 1630 3038
rect 1644 3036 1646 3038
rect 1649 3035 1651 3038
rect 1665 3036 1667 3038
rect 1681 3036 1683 3038
rect 1686 3033 1688 3038
rect 1707 3033 1709 3038
rect 1723 3036 1725 3038
rect 1739 3036 1741 3038
rect 1744 3033 1746 3038
rect 1760 3036 1762 3038
rect 1776 3036 1778 3038
rect 1781 3035 1783 3038
rect 1797 3036 1799 3038
rect 1813 3036 1815 3038
rect 1818 3033 1820 3038
rect 1839 3033 1841 3038
rect 1855 3036 1857 3038
rect 1871 3036 1873 3038
rect 1876 3033 1878 3038
rect 1892 3036 1894 3038
rect 2457 3036 2459 3038
rect 2462 3035 2464 3038
rect 2478 3036 2480 3038
rect 2494 3036 2496 3038
rect 2499 3033 2501 3038
rect 2520 3033 2522 3038
rect 2536 3036 2538 3038
rect 2552 3036 2554 3038
rect 2557 3033 2559 3038
rect 2573 3036 2575 3038
rect 2589 3036 2591 3038
rect 2594 3035 2596 3038
rect 2610 3036 2612 3038
rect 2626 3036 2628 3038
rect 2631 3033 2633 3038
rect 2652 3033 2654 3038
rect 2668 3036 2670 3038
rect 2684 3036 2686 3038
rect 2689 3033 2691 3038
rect 2705 3036 2707 3038
rect 2721 3036 2723 3038
rect 2726 3035 2728 3038
rect 2742 3036 2744 3038
rect 2758 3036 2760 3038
rect 2763 3033 2765 3038
rect 2784 3033 2786 3038
rect 2800 3036 2802 3038
rect 2816 3036 2818 3038
rect 2821 3033 2823 3038
rect 2837 3036 2839 3038
rect 2295 3013 2297 3015
rect 2300 3013 2302 3016
rect 2316 3013 2318 3015
rect 2332 3013 2334 3015
rect 2337 3013 2339 3016
rect 2358 3013 2360 3016
rect 2374 3013 2376 3016
rect 2390 3013 2392 3015
rect 2395 3013 2397 3016
rect 2411 3013 2413 3015
rect 3240 3013 3242 3015
rect 3245 3013 3247 3016
rect 3261 3013 3263 3015
rect 3277 3013 3279 3015
rect 3282 3013 3284 3016
rect 3303 3013 3305 3016
rect 3319 3013 3321 3016
rect 3335 3013 3337 3015
rect 3340 3013 3342 3016
rect 3356 3013 3358 3015
rect 2295 3000 2297 3005
rect 2300 3003 2302 3005
rect 2295 2986 2297 2996
rect 2300 2986 2302 2993
rect 2316 2986 2318 3005
rect 2332 2996 2334 3005
rect 2337 3003 2339 3005
rect 2358 3003 2360 3005
rect 2374 3002 2376 3005
rect 2332 2986 2334 2989
rect 2337 2986 2339 2988
rect 2358 2986 2360 2988
rect 2374 2986 2376 2998
rect 2390 2996 2392 3005
rect 2395 3003 2397 3005
rect 2390 2986 2392 2989
rect 2395 2986 2397 2988
rect 2411 2986 2413 3005
rect 3240 3000 3242 3005
rect 3245 3003 3247 3005
rect 2433 2992 2436 2994
rect 2440 2992 2443 2994
rect 3240 2986 3242 2996
rect 3245 2986 3247 2993
rect 3261 2986 3263 3005
rect 3277 2996 3279 3005
rect 3282 3003 3284 3005
rect 3303 3003 3305 3005
rect 3319 3002 3321 3005
rect 3277 2986 3279 2989
rect 3282 2986 3284 2988
rect 3303 2986 3305 2988
rect 3319 2986 3321 2998
rect 3335 2996 3337 3005
rect 3340 3003 3342 3005
rect 3335 2986 3337 2989
rect 3340 2986 3342 2988
rect 3356 2986 3358 3005
rect 3378 2992 3381 2994
rect 3385 2992 3388 2994
rect 1512 2983 1514 2985
rect 1517 2983 1519 2986
rect 1533 2983 1535 2985
rect 1549 2983 1551 2985
rect 1554 2983 1556 2986
rect 1575 2983 1577 2986
rect 1591 2983 1593 2986
rect 1607 2983 1609 2985
rect 1612 2983 1614 2986
rect 1628 2983 1630 2985
rect 1644 2983 1646 2985
rect 1649 2983 1651 2986
rect 1665 2983 1667 2985
rect 1681 2983 1683 2985
rect 1686 2983 1688 2986
rect 1707 2983 1709 2986
rect 1723 2983 1725 2986
rect 1739 2983 1741 2985
rect 1744 2983 1746 2986
rect 1760 2983 1762 2985
rect 1776 2983 1778 2985
rect 1781 2983 1783 2986
rect 1797 2983 1799 2985
rect 1813 2983 1815 2985
rect 1818 2983 1820 2986
rect 1839 2983 1841 2986
rect 1855 2983 1857 2986
rect 1871 2983 1873 2985
rect 1876 2983 1878 2986
rect 1892 2983 1894 2985
rect 2457 2983 2459 2985
rect 2462 2983 2464 2986
rect 2478 2983 2480 2985
rect 2494 2983 2496 2985
rect 2499 2983 2501 2986
rect 2520 2983 2522 2986
rect 2536 2983 2538 2986
rect 2552 2983 2554 2985
rect 2557 2983 2559 2986
rect 2573 2983 2575 2985
rect 2589 2983 2591 2985
rect 2594 2983 2596 2986
rect 2610 2983 2612 2985
rect 2626 2983 2628 2985
rect 2631 2983 2633 2986
rect 2652 2983 2654 2986
rect 2668 2983 2670 2986
rect 2684 2983 2686 2985
rect 2689 2983 2691 2986
rect 2705 2983 2707 2985
rect 2721 2983 2723 2985
rect 2726 2983 2728 2986
rect 2742 2983 2744 2985
rect 2758 2983 2760 2985
rect 2763 2983 2765 2986
rect 2784 2983 2786 2986
rect 2800 2983 2802 2986
rect 2816 2983 2818 2985
rect 2821 2983 2823 2986
rect 2837 2983 2839 2985
rect 2295 2980 2297 2982
rect 2300 2979 2302 2982
rect 2316 2980 2318 2982
rect 2332 2980 2334 2982
rect 2337 2977 2339 2982
rect 2358 2977 2360 2982
rect 2374 2980 2376 2982
rect 2390 2980 2392 2982
rect 2395 2977 2397 2982
rect 2411 2980 2413 2982
rect 1512 2970 1514 2975
rect 1517 2973 1519 2975
rect 1512 2956 1514 2966
rect 1517 2956 1519 2963
rect 1533 2956 1535 2975
rect 1549 2966 1551 2975
rect 1554 2973 1556 2975
rect 1575 2973 1577 2975
rect 1591 2972 1593 2975
rect 1549 2956 1551 2959
rect 1554 2956 1556 2958
rect 1575 2956 1577 2958
rect 1591 2956 1593 2968
rect 1607 2966 1609 2975
rect 1612 2973 1614 2975
rect 1607 2956 1609 2959
rect 1612 2956 1614 2958
rect 1628 2956 1630 2975
rect 1644 2972 1646 2975
rect 1649 2973 1651 2975
rect 1644 2956 1646 2968
rect 1649 2956 1651 2963
rect 1665 2956 1667 2975
rect 1681 2966 1683 2975
rect 1686 2973 1688 2975
rect 1707 2973 1709 2975
rect 1723 2972 1725 2975
rect 1681 2956 1683 2959
rect 1686 2956 1688 2958
rect 1707 2956 1709 2958
rect 1723 2956 1725 2968
rect 1739 2966 1741 2975
rect 1744 2973 1746 2975
rect 1739 2956 1741 2959
rect 1744 2956 1746 2958
rect 1760 2956 1762 2975
rect 1776 2972 1778 2975
rect 1781 2973 1783 2975
rect 1776 2956 1778 2968
rect 1781 2956 1783 2963
rect 1797 2956 1799 2975
rect 1813 2966 1815 2975
rect 1818 2973 1820 2975
rect 1839 2973 1841 2975
rect 1855 2972 1857 2975
rect 1813 2956 1815 2959
rect 1818 2956 1820 2958
rect 1839 2956 1841 2958
rect 1855 2956 1857 2968
rect 1871 2966 1873 2975
rect 1876 2973 1878 2975
rect 1892 2967 1894 2975
rect 3240 2980 3242 2982
rect 3245 2979 3247 2982
rect 3261 2980 3263 2982
rect 3277 2980 3279 2982
rect 3282 2977 3284 2982
rect 3303 2977 3305 2982
rect 3319 2980 3321 2982
rect 3335 2980 3337 2982
rect 3340 2977 3342 2982
rect 3356 2980 3358 2982
rect 2457 2970 2459 2975
rect 2462 2973 2464 2975
rect 1871 2956 1873 2959
rect 1876 2956 1878 2958
rect 1892 2956 1894 2963
rect 2457 2956 2459 2966
rect 2462 2956 2464 2963
rect 2478 2956 2480 2975
rect 2494 2966 2496 2975
rect 2499 2973 2501 2975
rect 2520 2973 2522 2975
rect 2536 2972 2538 2975
rect 2494 2956 2496 2959
rect 2499 2956 2501 2958
rect 2520 2956 2522 2958
rect 2536 2956 2538 2968
rect 2552 2966 2554 2975
rect 2557 2973 2559 2975
rect 2552 2956 2554 2959
rect 2557 2956 2559 2958
rect 2573 2956 2575 2975
rect 2589 2972 2591 2975
rect 2594 2973 2596 2975
rect 2589 2956 2591 2968
rect 2594 2956 2596 2963
rect 2610 2956 2612 2975
rect 2626 2966 2628 2975
rect 2631 2973 2633 2975
rect 2652 2973 2654 2975
rect 2668 2972 2670 2975
rect 2626 2956 2628 2959
rect 2631 2956 2633 2958
rect 2652 2956 2654 2958
rect 2668 2956 2670 2968
rect 2684 2966 2686 2975
rect 2689 2973 2691 2975
rect 2684 2956 2686 2959
rect 2689 2956 2691 2958
rect 2705 2956 2707 2975
rect 2721 2972 2723 2975
rect 2726 2973 2728 2975
rect 2721 2956 2723 2968
rect 2726 2956 2728 2963
rect 2742 2956 2744 2975
rect 2758 2966 2760 2975
rect 2763 2973 2765 2975
rect 2784 2973 2786 2975
rect 2800 2972 2802 2975
rect 2758 2956 2760 2959
rect 2763 2956 2765 2958
rect 2784 2956 2786 2958
rect 2800 2956 2802 2968
rect 2816 2966 2818 2975
rect 2821 2973 2823 2975
rect 2837 2967 2839 2975
rect 2816 2956 2818 2959
rect 2821 2956 2823 2958
rect 2837 2956 2839 2963
rect 1512 2950 1514 2952
rect 1517 2949 1519 2952
rect 1533 2950 1535 2952
rect 1549 2950 1551 2952
rect 1554 2947 1556 2952
rect 1575 2947 1577 2952
rect 1591 2950 1593 2952
rect 1607 2950 1609 2952
rect 1612 2947 1614 2952
rect 1628 2950 1630 2952
rect 1644 2950 1646 2952
rect 1649 2949 1651 2952
rect 1665 2950 1667 2952
rect 1681 2950 1683 2952
rect 1686 2947 1688 2952
rect 1707 2947 1709 2952
rect 1723 2950 1725 2952
rect 1739 2950 1741 2952
rect 1744 2947 1746 2952
rect 1760 2950 1762 2952
rect 1776 2950 1778 2952
rect 1781 2949 1783 2952
rect 1797 2950 1799 2952
rect 1813 2950 1815 2952
rect 1818 2947 1820 2952
rect 1839 2947 1841 2952
rect 1855 2950 1857 2952
rect 1871 2950 1873 2952
rect 1876 2947 1878 2952
rect 1892 2950 1894 2952
rect 2457 2950 2459 2952
rect 2462 2949 2464 2952
rect 2478 2950 2480 2952
rect 2494 2950 2496 2952
rect 2499 2947 2501 2952
rect 2520 2947 2522 2952
rect 2536 2950 2538 2952
rect 2552 2950 2554 2952
rect 2557 2947 2559 2952
rect 2573 2950 2575 2952
rect 2589 2950 2591 2952
rect 2594 2949 2596 2952
rect 2610 2950 2612 2952
rect 2626 2950 2628 2952
rect 2631 2947 2633 2952
rect 2652 2947 2654 2952
rect 2668 2950 2670 2952
rect 2684 2950 2686 2952
rect 2689 2947 2691 2952
rect 2705 2950 2707 2952
rect 2721 2950 2723 2952
rect 2726 2949 2728 2952
rect 2742 2950 2744 2952
rect 2758 2950 2760 2952
rect 2763 2947 2765 2952
rect 2784 2947 2786 2952
rect 2800 2950 2802 2952
rect 2816 2950 2818 2952
rect 2821 2947 2823 2952
rect 2837 2950 2839 2952
rect 1744 2912 1746 2915
rect 1768 2912 1770 2915
rect 2689 2912 2691 2915
rect 2713 2912 2715 2915
rect 1744 2906 1746 2908
rect 1768 2906 1770 2908
rect 2689 2906 2691 2908
rect 2713 2906 2715 2908
rect 1764 2901 1766 2903
rect 2709 2901 2711 2903
rect 1764 2894 1766 2897
rect 2709 2894 2711 2897
rect 1753 2883 1755 2885
rect 1759 2883 1778 2885
rect 2698 2883 2700 2885
rect 2704 2883 2723 2885
rect 1744 2878 1746 2880
rect 1768 2878 1770 2880
rect 2689 2878 2691 2880
rect 2713 2878 2715 2880
rect 1744 2871 1746 2874
rect 1768 2871 1770 2874
rect 2689 2871 2691 2874
rect 2713 2871 2715 2874
rect 1512 2843 1514 2845
rect 1517 2843 1519 2846
rect 1533 2843 1535 2845
rect 1549 2843 1551 2845
rect 1554 2843 1556 2846
rect 1575 2843 1577 2846
rect 1591 2843 1593 2846
rect 1607 2843 1609 2845
rect 1612 2843 1614 2846
rect 1628 2843 1630 2845
rect 1644 2843 1646 2845
rect 1649 2843 1651 2846
rect 1665 2843 1667 2845
rect 1681 2843 1683 2845
rect 1686 2843 1688 2846
rect 1707 2843 1709 2846
rect 1723 2843 1725 2846
rect 1739 2843 1741 2845
rect 1744 2843 1746 2846
rect 1760 2843 1762 2845
rect 1776 2843 1778 2845
rect 1781 2843 1783 2846
rect 1797 2843 1799 2845
rect 1813 2843 1815 2845
rect 1818 2843 1820 2846
rect 1839 2843 1841 2846
rect 1855 2843 1857 2846
rect 1871 2843 1873 2845
rect 1876 2843 1878 2846
rect 1892 2843 1894 2845
rect 2457 2843 2459 2845
rect 2462 2843 2464 2846
rect 2478 2843 2480 2845
rect 2494 2843 2496 2845
rect 2499 2843 2501 2846
rect 2520 2843 2522 2846
rect 2536 2843 2538 2846
rect 2552 2843 2554 2845
rect 2557 2843 2559 2846
rect 2573 2843 2575 2845
rect 2589 2843 2591 2845
rect 2594 2843 2596 2846
rect 2610 2843 2612 2845
rect 2626 2843 2628 2845
rect 2631 2843 2633 2846
rect 2652 2843 2654 2846
rect 2668 2843 2670 2846
rect 2684 2843 2686 2845
rect 2689 2843 2691 2846
rect 2705 2843 2707 2845
rect 2721 2843 2723 2845
rect 2726 2843 2728 2846
rect 2742 2843 2744 2845
rect 2758 2843 2760 2845
rect 2763 2843 2765 2846
rect 2784 2843 2786 2846
rect 2800 2843 2802 2846
rect 2816 2843 2818 2845
rect 2821 2843 2823 2846
rect 2837 2843 2839 2845
rect 1512 2830 1514 2835
rect 1517 2833 1519 2835
rect 1512 2816 1514 2826
rect 1517 2816 1519 2823
rect 1533 2816 1535 2835
rect 1549 2826 1551 2835
rect 1554 2833 1556 2835
rect 1575 2833 1577 2835
rect 1591 2832 1593 2835
rect 1549 2816 1551 2819
rect 1554 2816 1556 2818
rect 1575 2816 1577 2818
rect 1591 2816 1593 2828
rect 1607 2826 1609 2835
rect 1612 2833 1614 2835
rect 1607 2816 1609 2819
rect 1612 2816 1614 2818
rect 1628 2816 1630 2835
rect 1644 2832 1646 2835
rect 1649 2833 1651 2835
rect 1644 2816 1646 2828
rect 1649 2816 1651 2823
rect 1665 2816 1667 2835
rect 1681 2826 1683 2835
rect 1686 2833 1688 2835
rect 1707 2833 1709 2835
rect 1723 2832 1725 2835
rect 1681 2816 1683 2819
rect 1686 2816 1688 2818
rect 1707 2816 1709 2818
rect 1723 2816 1725 2828
rect 1739 2826 1741 2835
rect 1744 2833 1746 2835
rect 1739 2816 1741 2819
rect 1744 2816 1746 2818
rect 1760 2816 1762 2835
rect 1776 2832 1778 2835
rect 1781 2833 1783 2835
rect 1776 2816 1778 2828
rect 1781 2816 1783 2823
rect 1797 2816 1799 2835
rect 1813 2826 1815 2835
rect 1818 2833 1820 2835
rect 1839 2833 1841 2835
rect 1855 2832 1857 2835
rect 1813 2816 1815 2819
rect 1818 2816 1820 2818
rect 1839 2816 1841 2818
rect 1855 2816 1857 2828
rect 1871 2826 1873 2835
rect 1876 2833 1878 2835
rect 1892 2827 1894 2835
rect 2457 2830 2459 2835
rect 2462 2833 2464 2835
rect 1871 2816 1873 2819
rect 1876 2816 1878 2818
rect 1892 2816 1894 2823
rect 2457 2816 2459 2826
rect 2462 2816 2464 2823
rect 2478 2816 2480 2835
rect 2494 2826 2496 2835
rect 2499 2833 2501 2835
rect 2520 2833 2522 2835
rect 2536 2832 2538 2835
rect 2494 2816 2496 2819
rect 2499 2816 2501 2818
rect 2520 2816 2522 2818
rect 2536 2816 2538 2828
rect 2552 2826 2554 2835
rect 2557 2833 2559 2835
rect 2552 2816 2554 2819
rect 2557 2816 2559 2818
rect 2573 2816 2575 2835
rect 2589 2832 2591 2835
rect 2594 2833 2596 2835
rect 2589 2816 2591 2828
rect 2594 2816 2596 2823
rect 2610 2816 2612 2835
rect 2626 2826 2628 2835
rect 2631 2833 2633 2835
rect 2652 2833 2654 2835
rect 2668 2832 2670 2835
rect 2626 2816 2628 2819
rect 2631 2816 2633 2818
rect 2652 2816 2654 2818
rect 2668 2816 2670 2828
rect 2684 2826 2686 2835
rect 2689 2833 2691 2835
rect 2684 2816 2686 2819
rect 2689 2816 2691 2818
rect 2705 2816 2707 2835
rect 2721 2832 2723 2835
rect 2726 2833 2728 2835
rect 2721 2816 2723 2828
rect 2726 2816 2728 2823
rect 2742 2816 2744 2835
rect 2758 2826 2760 2835
rect 2763 2833 2765 2835
rect 2784 2833 2786 2835
rect 2800 2832 2802 2835
rect 2758 2816 2760 2819
rect 2763 2816 2765 2818
rect 2784 2816 2786 2818
rect 2800 2816 2802 2828
rect 2816 2826 2818 2835
rect 2821 2833 2823 2835
rect 2837 2827 2839 2835
rect 2816 2816 2818 2819
rect 2821 2816 2823 2818
rect 2837 2816 2839 2823
rect 1512 2810 1514 2812
rect 1517 2809 1519 2812
rect 1533 2810 1535 2812
rect 1549 2810 1551 2812
rect 1554 2807 1556 2812
rect 1575 2807 1577 2812
rect 1591 2810 1593 2812
rect 1607 2810 1609 2812
rect 1612 2807 1614 2812
rect 1628 2810 1630 2812
rect 1644 2810 1646 2812
rect 1649 2809 1651 2812
rect 1665 2810 1667 2812
rect 1681 2810 1683 2812
rect 1686 2807 1688 2812
rect 1707 2807 1709 2812
rect 1723 2810 1725 2812
rect 1739 2810 1741 2812
rect 1744 2807 1746 2812
rect 1760 2810 1762 2812
rect 1776 2810 1778 2812
rect 1781 2809 1783 2812
rect 1797 2810 1799 2812
rect 1813 2810 1815 2812
rect 1818 2807 1820 2812
rect 1839 2807 1841 2812
rect 1855 2810 1857 2812
rect 1871 2810 1873 2812
rect 1876 2807 1878 2812
rect 1892 2810 1894 2812
rect 2457 2810 2459 2812
rect 2462 2809 2464 2812
rect 2478 2810 2480 2812
rect 2494 2810 2496 2812
rect 2499 2807 2501 2812
rect 2520 2807 2522 2812
rect 2536 2810 2538 2812
rect 2552 2810 2554 2812
rect 2557 2807 2559 2812
rect 2573 2810 2575 2812
rect 2589 2810 2591 2812
rect 2594 2809 2596 2812
rect 2610 2810 2612 2812
rect 2626 2810 2628 2812
rect 2631 2807 2633 2812
rect 2652 2807 2654 2812
rect 2668 2810 2670 2812
rect 2684 2810 2686 2812
rect 2689 2807 2691 2812
rect 2705 2810 2707 2812
rect 2721 2810 2723 2812
rect 2726 2809 2728 2812
rect 2742 2810 2744 2812
rect 2758 2810 2760 2812
rect 2763 2807 2765 2812
rect 2784 2807 2786 2812
rect 2800 2810 2802 2812
rect 2816 2810 2818 2812
rect 2821 2807 2823 2812
rect 2837 2810 2839 2812
rect 1996 2764 1998 2766
rect 2001 2764 2003 2767
rect 2017 2764 2019 2766
rect 2033 2764 2035 2766
rect 2038 2764 2040 2767
rect 2059 2764 2061 2767
rect 2075 2764 2077 2767
rect 2091 2764 2093 2766
rect 2096 2764 2098 2767
rect 2112 2764 2114 2766
rect 2128 2764 2130 2766
rect 2133 2764 2135 2767
rect 2149 2764 2151 2766
rect 2165 2764 2167 2766
rect 2170 2764 2172 2767
rect 2191 2764 2193 2767
rect 2207 2764 2209 2767
rect 2223 2764 2225 2766
rect 2228 2764 2230 2767
rect 2244 2764 2246 2766
rect 2260 2764 2262 2766
rect 2265 2764 2267 2767
rect 2281 2764 2283 2766
rect 2297 2764 2299 2766
rect 2302 2764 2304 2767
rect 2323 2764 2325 2767
rect 2339 2764 2341 2767
rect 2355 2764 2357 2766
rect 2360 2764 2362 2767
rect 2376 2764 2378 2766
rect 2392 2764 2394 2766
rect 2397 2764 2399 2767
rect 2413 2764 2415 2766
rect 2429 2764 2431 2766
rect 2434 2764 2436 2767
rect 2455 2764 2457 2767
rect 2471 2764 2473 2767
rect 2487 2764 2489 2766
rect 2492 2764 2494 2767
rect 2508 2764 2510 2766
rect 2941 2764 2943 2766
rect 2946 2764 2948 2767
rect 2962 2764 2964 2766
rect 2978 2764 2980 2766
rect 2983 2764 2985 2767
rect 3004 2764 3006 2767
rect 3020 2764 3022 2767
rect 3036 2764 3038 2766
rect 3041 2764 3043 2767
rect 3057 2764 3059 2766
rect 3073 2764 3075 2766
rect 3078 2764 3080 2767
rect 3094 2764 3096 2766
rect 3110 2764 3112 2766
rect 3115 2764 3117 2767
rect 3136 2764 3138 2767
rect 3152 2764 3154 2767
rect 3168 2764 3170 2766
rect 3173 2764 3175 2767
rect 3189 2764 3191 2766
rect 3205 2764 3207 2766
rect 3210 2764 3212 2767
rect 3226 2764 3228 2766
rect 3242 2764 3244 2766
rect 3247 2764 3249 2767
rect 3268 2764 3270 2767
rect 3284 2764 3286 2767
rect 3300 2764 3302 2766
rect 3305 2764 3307 2767
rect 3321 2764 3323 2766
rect 3337 2764 3339 2766
rect 3342 2764 3344 2767
rect 3358 2764 3360 2766
rect 3374 2764 3376 2766
rect 3379 2764 3381 2767
rect 3400 2764 3402 2767
rect 3416 2764 3418 2767
rect 3432 2764 3434 2766
rect 3437 2764 3439 2767
rect 3453 2764 3455 2766
rect 1996 2751 1998 2756
rect 2001 2754 2003 2756
rect 1996 2737 1998 2747
rect 2001 2737 2003 2744
rect 2017 2737 2019 2756
rect 2033 2747 2035 2756
rect 2038 2754 2040 2756
rect 2059 2754 2061 2756
rect 2075 2753 2077 2756
rect 2033 2737 2035 2740
rect 2038 2737 2040 2739
rect 2059 2737 2061 2739
rect 2075 2737 2077 2749
rect 2091 2747 2093 2756
rect 2096 2754 2098 2756
rect 2112 2748 2114 2756
rect 2128 2751 2130 2756
rect 2133 2754 2135 2756
rect 2091 2737 2093 2740
rect 2096 2737 2098 2739
rect 2112 2737 2114 2744
rect 2128 2737 2130 2747
rect 2133 2737 2135 2744
rect 2149 2737 2151 2756
rect 2165 2747 2167 2756
rect 2170 2754 2172 2756
rect 2191 2754 2193 2756
rect 2207 2753 2209 2756
rect 2165 2737 2167 2740
rect 2170 2737 2172 2739
rect 2191 2737 2193 2739
rect 2207 2737 2209 2749
rect 2223 2747 2225 2756
rect 2228 2754 2230 2756
rect 2244 2748 2246 2756
rect 2260 2751 2262 2756
rect 2265 2754 2267 2756
rect 2223 2737 2225 2740
rect 2228 2737 2230 2739
rect 2244 2737 2246 2744
rect 2260 2737 2262 2747
rect 2265 2737 2267 2744
rect 2281 2737 2283 2756
rect 2297 2747 2299 2756
rect 2302 2754 2304 2756
rect 2323 2754 2325 2756
rect 2339 2753 2341 2756
rect 2297 2737 2299 2740
rect 2302 2737 2304 2739
rect 2323 2737 2325 2739
rect 2339 2737 2341 2749
rect 2355 2747 2357 2756
rect 2360 2754 2362 2756
rect 2376 2748 2378 2756
rect 2392 2751 2394 2756
rect 2397 2754 2399 2756
rect 2355 2737 2357 2740
rect 2360 2737 2362 2739
rect 2376 2737 2378 2744
rect 2392 2737 2394 2747
rect 2397 2737 2399 2744
rect 2413 2737 2415 2756
rect 2429 2747 2431 2756
rect 2434 2754 2436 2756
rect 2455 2754 2457 2756
rect 2471 2753 2473 2756
rect 2429 2737 2431 2740
rect 2434 2737 2436 2739
rect 2455 2737 2457 2739
rect 2471 2737 2473 2749
rect 2487 2747 2489 2756
rect 2492 2754 2494 2756
rect 2508 2748 2510 2756
rect 2941 2751 2943 2756
rect 2946 2754 2948 2756
rect 2487 2737 2489 2740
rect 2492 2737 2494 2739
rect 2508 2737 2510 2744
rect 1644 2731 1646 2733
rect 1649 2731 1651 2734
rect 1665 2731 1667 2733
rect 1681 2731 1683 2733
rect 1686 2731 1688 2734
rect 1707 2731 1709 2734
rect 1723 2731 1725 2734
rect 1739 2731 1741 2733
rect 1744 2731 1746 2734
rect 2941 2737 2943 2747
rect 2946 2737 2948 2744
rect 2962 2737 2964 2756
rect 2978 2747 2980 2756
rect 2983 2754 2985 2756
rect 3004 2754 3006 2756
rect 3020 2753 3022 2756
rect 2978 2737 2980 2740
rect 2983 2737 2985 2739
rect 3004 2737 3006 2739
rect 3020 2737 3022 2749
rect 3036 2747 3038 2756
rect 3041 2754 3043 2756
rect 3057 2748 3059 2756
rect 3073 2751 3075 2756
rect 3078 2754 3080 2756
rect 3036 2737 3038 2740
rect 3041 2737 3043 2739
rect 3057 2737 3059 2744
rect 3073 2737 3075 2747
rect 3078 2737 3080 2744
rect 3094 2737 3096 2756
rect 3110 2747 3112 2756
rect 3115 2754 3117 2756
rect 3136 2754 3138 2756
rect 3152 2753 3154 2756
rect 3110 2737 3112 2740
rect 3115 2737 3117 2739
rect 3136 2737 3138 2739
rect 3152 2737 3154 2749
rect 3168 2747 3170 2756
rect 3173 2754 3175 2756
rect 3189 2748 3191 2756
rect 3205 2751 3207 2756
rect 3210 2754 3212 2756
rect 3168 2737 3170 2740
rect 3173 2737 3175 2739
rect 3189 2737 3191 2744
rect 3205 2737 3207 2747
rect 3210 2737 3212 2744
rect 3226 2737 3228 2756
rect 3242 2747 3244 2756
rect 3247 2754 3249 2756
rect 3268 2754 3270 2756
rect 3284 2753 3286 2756
rect 3242 2737 3244 2740
rect 3247 2737 3249 2739
rect 3268 2737 3270 2739
rect 3284 2737 3286 2749
rect 3300 2747 3302 2756
rect 3305 2754 3307 2756
rect 3321 2748 3323 2756
rect 3337 2751 3339 2756
rect 3342 2754 3344 2756
rect 3300 2737 3302 2740
rect 3305 2737 3307 2739
rect 3321 2737 3323 2744
rect 3337 2737 3339 2747
rect 3342 2737 3344 2744
rect 3358 2737 3360 2756
rect 3374 2747 3376 2756
rect 3379 2754 3381 2756
rect 3400 2754 3402 2756
rect 3416 2753 3418 2756
rect 3374 2737 3376 2740
rect 3379 2737 3381 2739
rect 3400 2737 3402 2739
rect 3416 2737 3418 2749
rect 3432 2747 3434 2756
rect 3437 2754 3439 2756
rect 3453 2748 3455 2756
rect 3432 2737 3434 2740
rect 3437 2737 3439 2739
rect 3453 2737 3455 2744
rect 1760 2731 1762 2733
rect 1996 2731 1998 2733
rect 2001 2730 2003 2733
rect 2017 2731 2019 2733
rect 2033 2731 2035 2733
rect 2038 2728 2040 2733
rect 2059 2728 2061 2733
rect 2075 2731 2077 2733
rect 2091 2731 2093 2733
rect 2096 2728 2098 2733
rect 2112 2731 2114 2733
rect 2128 2731 2130 2733
rect 2133 2730 2135 2733
rect 2149 2731 2151 2733
rect 2165 2731 2167 2733
rect 2170 2728 2172 2733
rect 2191 2728 2193 2733
rect 2207 2731 2209 2733
rect 2223 2731 2225 2733
rect 2228 2728 2230 2733
rect 2244 2731 2246 2733
rect 2260 2731 2262 2733
rect 2265 2730 2267 2733
rect 2281 2731 2283 2733
rect 2297 2731 2299 2733
rect 2302 2728 2304 2733
rect 2323 2728 2325 2733
rect 2339 2731 2341 2733
rect 2355 2731 2357 2733
rect 2360 2728 2362 2733
rect 2376 2731 2378 2733
rect 2392 2731 2394 2733
rect 2397 2730 2399 2733
rect 2413 2731 2415 2733
rect 2429 2731 2431 2733
rect 2434 2728 2436 2733
rect 2455 2728 2457 2733
rect 2471 2731 2473 2733
rect 2487 2731 2489 2733
rect 2492 2728 2494 2733
rect 2508 2731 2510 2733
rect 2589 2731 2591 2733
rect 2594 2731 2596 2734
rect 2610 2731 2612 2733
rect 2626 2731 2628 2733
rect 2631 2731 2633 2734
rect 2652 2731 2654 2734
rect 2668 2731 2670 2734
rect 2684 2731 2686 2733
rect 2689 2731 2691 2734
rect 2705 2731 2707 2733
rect 2941 2731 2943 2733
rect 2946 2730 2948 2733
rect 2962 2731 2964 2733
rect 2978 2731 2980 2733
rect 2983 2728 2985 2733
rect 3004 2728 3006 2733
rect 3020 2731 3022 2733
rect 3036 2731 3038 2733
rect 3041 2728 3043 2733
rect 3057 2731 3059 2733
rect 3073 2731 3075 2733
rect 3078 2730 3080 2733
rect 3094 2731 3096 2733
rect 3110 2731 3112 2733
rect 3115 2728 3117 2733
rect 3136 2728 3138 2733
rect 3152 2731 3154 2733
rect 3168 2731 3170 2733
rect 3173 2728 3175 2733
rect 3189 2731 3191 2733
rect 3205 2731 3207 2733
rect 3210 2730 3212 2733
rect 3226 2731 3228 2733
rect 3242 2731 3244 2733
rect 3247 2728 3249 2733
rect 3268 2728 3270 2733
rect 3284 2731 3286 2733
rect 3300 2731 3302 2733
rect 3305 2728 3307 2733
rect 3321 2731 3323 2733
rect 3337 2731 3339 2733
rect 3342 2730 3344 2733
rect 3358 2731 3360 2733
rect 3374 2731 3376 2733
rect 3379 2728 3381 2733
rect 3400 2728 3402 2733
rect 3416 2731 3418 2733
rect 3432 2731 3434 2733
rect 3437 2728 3439 2733
rect 3453 2731 3455 2733
rect 1644 2718 1646 2723
rect 1649 2721 1651 2723
rect 1644 2704 1646 2714
rect 1649 2704 1651 2711
rect 1665 2704 1667 2723
rect 1681 2714 1683 2723
rect 1686 2721 1688 2723
rect 1707 2721 1709 2723
rect 1723 2720 1725 2723
rect 1681 2704 1683 2707
rect 1686 2704 1688 2706
rect 1707 2704 1709 2706
rect 1723 2704 1725 2716
rect 1739 2714 1741 2723
rect 1744 2721 1746 2723
rect 1739 2704 1741 2707
rect 1744 2704 1746 2706
rect 1760 2704 1762 2723
rect 2589 2718 2591 2723
rect 2594 2721 2596 2723
rect 2589 2704 2591 2714
rect 2594 2704 2596 2711
rect 2610 2704 2612 2723
rect 2626 2714 2628 2723
rect 2631 2721 2633 2723
rect 2652 2721 2654 2723
rect 2668 2720 2670 2723
rect 2626 2704 2628 2707
rect 2631 2704 2633 2706
rect 2652 2704 2654 2706
rect 2668 2704 2670 2716
rect 2684 2714 2686 2723
rect 2689 2721 2691 2723
rect 2684 2704 2686 2707
rect 2689 2704 2691 2706
rect 2705 2704 2707 2723
rect 1644 2698 1646 2700
rect 1649 2697 1651 2700
rect 1665 2698 1667 2700
rect 1681 2698 1683 2700
rect 1686 2695 1688 2700
rect 1707 2695 1709 2700
rect 1723 2698 1725 2700
rect 1739 2698 1741 2700
rect 1744 2695 1746 2700
rect 1760 2698 1762 2700
rect 2589 2698 2591 2700
rect 2594 2697 2596 2700
rect 2610 2698 2612 2700
rect 2626 2698 2628 2700
rect 2175 2693 2177 2695
rect 2017 2687 2019 2690
rect 2061 2687 2063 2690
rect 2087 2687 2089 2690
rect 2133 2687 2135 2690
rect 2087 2683 2088 2687
rect 2201 2687 2203 2691
rect 2229 2693 2231 2695
rect 2256 2693 2258 2695
rect 2206 2687 2208 2690
rect 2001 2680 2003 2682
rect 2017 2680 2019 2683
rect 2033 2680 2035 2682
rect 2056 2680 2058 2682
rect 2061 2680 2063 2683
rect 2087 2680 2089 2683
rect 2108 2680 2110 2683
rect 2128 2680 2130 2682
rect 2133 2680 2135 2683
rect 2151 2680 2153 2682
rect 1768 2667 1770 2670
rect 1768 2661 1770 2663
rect 1651 2658 1653 2661
rect 2001 2658 2003 2672
rect 2017 2670 2019 2672
rect 2017 2658 2019 2660
rect 2033 2658 2035 2672
rect 2056 2667 2058 2672
rect 2061 2670 2063 2672
rect 2087 2670 2089 2672
rect 2052 2663 2058 2667
rect 2056 2658 2058 2663
rect 2061 2658 2063 2660
rect 2087 2658 2089 2660
rect 2108 2658 2110 2672
rect 2128 2667 2130 2672
rect 2133 2670 2135 2672
rect 2124 2663 2130 2667
rect 2128 2658 2130 2663
rect 2133 2658 2135 2660
rect 2151 2658 2153 2672
rect 2175 2671 2177 2685
rect 2282 2687 2284 2691
rect 2310 2693 2312 2695
rect 2631 2695 2633 2700
rect 2652 2695 2654 2700
rect 2668 2698 2670 2700
rect 2684 2698 2686 2700
rect 2689 2695 2691 2700
rect 2705 2698 2707 2700
rect 2287 2687 2289 2690
rect 2201 2676 2203 2679
rect 2206 2677 2208 2679
rect 2202 2672 2203 2676
rect 2201 2667 2203 2672
rect 2206 2667 2208 2669
rect 2175 2665 2177 2667
rect 2229 2663 2231 2685
rect 2256 2671 2258 2685
rect 3120 2693 3122 2695
rect 2282 2676 2284 2679
rect 2287 2677 2289 2679
rect 2283 2672 2284 2676
rect 2282 2667 2284 2672
rect 2287 2667 2289 2669
rect 2256 2665 2258 2667
rect 2310 2663 2312 2685
rect 2962 2687 2964 2690
rect 3006 2687 3008 2690
rect 3032 2687 3034 2690
rect 3078 2687 3080 2690
rect 3032 2683 3033 2687
rect 3146 2687 3148 2691
rect 3174 2693 3176 2695
rect 3201 2693 3203 2695
rect 3151 2687 3153 2690
rect 2946 2680 2948 2682
rect 2962 2680 2964 2683
rect 2978 2680 2980 2682
rect 3001 2680 3003 2682
rect 3006 2680 3008 2683
rect 3032 2680 3034 2683
rect 3053 2680 3055 2683
rect 3073 2680 3075 2682
rect 3078 2680 3080 2683
rect 3096 2680 3098 2682
rect 2713 2667 2715 2670
rect 2201 2661 2203 2663
rect 2206 2658 2208 2663
rect 2282 2661 2284 2663
rect 2229 2657 2231 2659
rect 2287 2658 2289 2663
rect 2713 2661 2715 2663
rect 2310 2657 2312 2659
rect 2596 2658 2598 2661
rect 2946 2658 2948 2672
rect 2962 2670 2964 2672
rect 2962 2658 2964 2660
rect 2978 2658 2980 2672
rect 3001 2667 3003 2672
rect 3006 2670 3008 2672
rect 3032 2670 3034 2672
rect 2997 2663 3003 2667
rect 3001 2658 3003 2663
rect 3006 2658 3008 2660
rect 3032 2658 3034 2660
rect 3053 2658 3055 2672
rect 3073 2667 3075 2672
rect 3078 2670 3080 2672
rect 3069 2663 3075 2667
rect 3073 2658 3075 2663
rect 3078 2658 3080 2660
rect 3096 2658 3098 2672
rect 3120 2671 3122 2685
rect 3227 2687 3229 2691
rect 3255 2693 3257 2695
rect 3232 2687 3234 2690
rect 3146 2676 3148 2679
rect 3151 2677 3153 2679
rect 3147 2672 3148 2676
rect 3146 2667 3148 2672
rect 3151 2667 3153 2669
rect 3120 2665 3122 2667
rect 3174 2663 3176 2685
rect 3201 2671 3203 2685
rect 3227 2676 3229 2679
rect 3232 2677 3234 2679
rect 3228 2672 3229 2676
rect 3227 2667 3229 2672
rect 3232 2667 3234 2669
rect 3201 2665 3203 2667
rect 3255 2663 3257 2685
rect 3146 2661 3148 2663
rect 3151 2658 3153 2663
rect 3227 2661 3229 2663
rect 3174 2657 3176 2659
rect 3232 2658 3234 2663
rect 3255 2657 3257 2659
rect 1651 2652 1653 2654
rect 2001 2652 2003 2654
rect 2017 2650 2019 2654
rect 2033 2652 2035 2654
rect 2056 2652 2058 2654
rect 2018 2646 2019 2650
rect 2061 2649 2063 2654
rect 2087 2650 2089 2654
rect 2108 2652 2110 2654
rect 2128 2652 2130 2654
rect 2017 2643 2019 2646
rect 2062 2645 2063 2649
rect 2088 2646 2089 2650
rect 2133 2649 2135 2654
rect 2151 2652 2153 2654
rect 2596 2652 2598 2654
rect 2946 2652 2948 2654
rect 2962 2650 2964 2654
rect 2978 2652 2980 2654
rect 3001 2652 3003 2654
rect 2061 2643 2063 2645
rect 2087 2642 2089 2646
rect 2134 2645 2135 2649
rect 2963 2646 2964 2650
rect 3006 2649 3008 2654
rect 3032 2650 3034 2654
rect 3053 2652 3055 2654
rect 3073 2652 3075 2654
rect 2133 2643 2135 2645
rect 2962 2643 2964 2646
rect 3007 2645 3008 2649
rect 3033 2646 3034 2650
rect 3078 2649 3080 2654
rect 3096 2652 3098 2654
rect 3006 2643 3008 2645
rect 3032 2642 3034 2646
rect 3079 2645 3080 2649
rect 3078 2643 3080 2645
rect 1635 2629 1637 2631
rect 1651 2629 1653 2632
rect 1656 2629 1658 2631
rect 1672 2629 1674 2632
rect 1688 2629 1690 2632
rect 1709 2629 1711 2632
rect 1714 2629 1716 2631
rect 1730 2629 1732 2631
rect 1746 2629 1748 2632
rect 1751 2629 1753 2631
rect 2580 2629 2582 2631
rect 2596 2629 2598 2632
rect 2601 2629 2603 2631
rect 2617 2629 2619 2632
rect 2633 2629 2635 2632
rect 2654 2629 2656 2632
rect 2659 2629 2661 2631
rect 2675 2629 2677 2631
rect 2691 2629 2693 2632
rect 2696 2629 2698 2631
rect 1635 2602 1637 2621
rect 1651 2619 1653 2621
rect 1656 2612 1658 2621
rect 1672 2618 1674 2621
rect 1688 2619 1690 2621
rect 1709 2619 1711 2621
rect 1651 2602 1653 2604
rect 1656 2602 1658 2605
rect 1672 2602 1674 2614
rect 1714 2612 1716 2621
rect 1688 2602 1690 2604
rect 1709 2602 1711 2604
rect 1714 2602 1716 2605
rect 1730 2602 1732 2621
rect 1746 2619 1748 2621
rect 1751 2616 1753 2621
rect 2017 2620 2019 2623
rect 2061 2621 2063 2623
rect 2018 2616 2019 2620
rect 2062 2617 2063 2621
rect 2087 2620 2089 2624
rect 2133 2621 2135 2623
rect 2001 2612 2003 2614
rect 2017 2612 2019 2616
rect 2033 2612 2035 2614
rect 2056 2612 2058 2614
rect 2061 2612 2063 2617
rect 2088 2616 2089 2620
rect 2134 2617 2135 2621
rect 2087 2612 2089 2616
rect 2108 2612 2110 2614
rect 2128 2612 2130 2614
rect 2133 2612 2135 2617
rect 2151 2612 2153 2614
rect 1746 2602 1748 2609
rect 1751 2602 1753 2612
rect 2201 2611 2203 2614
rect 2206 2611 2208 2614
rect 2282 2611 2284 2614
rect 2287 2611 2289 2614
rect 1635 2596 1637 2598
rect 1651 2593 1653 2598
rect 1656 2596 1658 2598
rect 1672 2596 1674 2598
rect 1688 2593 1690 2598
rect 1709 2593 1711 2598
rect 1714 2596 1716 2598
rect 1730 2596 1732 2598
rect 1746 2595 1748 2598
rect 1751 2596 1753 2598
rect 2001 2594 2003 2608
rect 2017 2606 2019 2608
rect 2017 2594 2019 2596
rect 2033 2594 2035 2608
rect 2056 2603 2058 2608
rect 2061 2606 2063 2608
rect 2087 2606 2089 2608
rect 2052 2599 2058 2603
rect 2056 2594 2058 2599
rect 2061 2594 2063 2596
rect 2087 2594 2089 2596
rect 2108 2594 2110 2608
rect 2128 2603 2130 2608
rect 2133 2606 2135 2608
rect 2124 2599 2130 2603
rect 2128 2594 2130 2599
rect 2133 2594 2135 2596
rect 2151 2594 2153 2608
rect 2201 2595 2203 2607
rect 2206 2605 2208 2607
rect 2206 2595 2208 2597
rect 2282 2595 2284 2607
rect 2287 2605 2289 2607
rect 2580 2602 2582 2621
rect 2596 2619 2598 2621
rect 2601 2612 2603 2621
rect 2617 2618 2619 2621
rect 2633 2619 2635 2621
rect 2654 2619 2656 2621
rect 2596 2602 2598 2604
rect 2601 2602 2603 2605
rect 2617 2602 2619 2614
rect 2659 2612 2661 2621
rect 2633 2602 2635 2604
rect 2654 2602 2656 2604
rect 2659 2602 2661 2605
rect 2675 2602 2677 2621
rect 2691 2619 2693 2621
rect 2696 2616 2698 2621
rect 2962 2620 2964 2623
rect 3006 2621 3008 2623
rect 2963 2616 2964 2620
rect 3007 2617 3008 2621
rect 3032 2620 3034 2624
rect 3078 2621 3080 2623
rect 2946 2612 2948 2614
rect 2962 2612 2964 2616
rect 2978 2612 2980 2614
rect 3001 2612 3003 2614
rect 3006 2612 3008 2617
rect 3033 2616 3034 2620
rect 3079 2617 3080 2621
rect 3032 2612 3034 2616
rect 3053 2612 3055 2614
rect 3073 2612 3075 2614
rect 3078 2612 3080 2617
rect 3096 2612 3098 2614
rect 2691 2602 2693 2609
rect 2696 2602 2698 2612
rect 3146 2611 3148 2614
rect 3151 2611 3153 2614
rect 3227 2611 3229 2614
rect 3232 2611 3234 2614
rect 2287 2595 2289 2597
rect 2580 2596 2582 2598
rect 2596 2593 2598 2598
rect 2601 2596 2603 2598
rect 2617 2596 2619 2598
rect 2633 2593 2635 2598
rect 2654 2593 2656 2598
rect 2659 2596 2661 2598
rect 2675 2596 2677 2598
rect 2691 2595 2693 2598
rect 2696 2596 2698 2598
rect 2946 2594 2948 2608
rect 2962 2606 2964 2608
rect 2962 2594 2964 2596
rect 2978 2594 2980 2608
rect 3001 2603 3003 2608
rect 3006 2606 3008 2608
rect 3032 2606 3034 2608
rect 2997 2599 3003 2603
rect 3001 2594 3003 2599
rect 3006 2594 3008 2596
rect 3032 2594 3034 2596
rect 3053 2594 3055 2608
rect 3073 2603 3075 2608
rect 3078 2606 3080 2608
rect 3069 2599 3075 2603
rect 3073 2594 3075 2599
rect 3078 2594 3080 2596
rect 3096 2594 3098 2608
rect 3146 2595 3148 2607
rect 3151 2605 3153 2607
rect 3151 2595 3153 2597
rect 3227 2595 3229 2607
rect 3232 2605 3234 2607
rect 3232 2595 3234 2597
rect 2001 2584 2003 2586
rect 2017 2583 2019 2586
rect 2033 2584 2035 2586
rect 2056 2584 2058 2586
rect 2061 2583 2063 2586
rect 2087 2583 2089 2586
rect 2108 2583 2110 2586
rect 2128 2584 2130 2586
rect 2133 2583 2135 2586
rect 2151 2584 2153 2586
rect 2201 2585 2203 2587
rect 2087 2579 2088 2583
rect 2206 2582 2208 2587
rect 2282 2585 2284 2587
rect 2287 2582 2289 2587
rect 2946 2584 2948 2586
rect 2962 2583 2964 2586
rect 2978 2584 2980 2586
rect 3001 2584 3003 2586
rect 3006 2583 3008 2586
rect 3032 2583 3034 2586
rect 3053 2583 3055 2586
rect 3073 2584 3075 2586
rect 3078 2583 3080 2586
rect 3096 2584 3098 2586
rect 3146 2585 3148 2587
rect 2017 2576 2019 2579
rect 2061 2576 2063 2579
rect 2087 2576 2089 2579
rect 2133 2576 2135 2579
rect 3032 2579 3033 2583
rect 3151 2582 3153 2587
rect 3227 2585 3229 2587
rect 3232 2582 3234 2587
rect 2962 2576 2964 2579
rect 3006 2576 3008 2579
rect 3032 2576 3034 2579
rect 3078 2576 3080 2579
rect 2017 2555 2019 2558
rect 2061 2555 2063 2558
rect 2087 2555 2089 2558
rect 2133 2555 2135 2558
rect 2201 2555 2203 2559
rect 2229 2561 2231 2563
rect 2280 2561 2282 2563
rect 2206 2555 2208 2558
rect 2087 2551 2088 2555
rect 2001 2548 2003 2550
rect 2017 2548 2019 2551
rect 2033 2548 2035 2550
rect 2056 2548 2058 2550
rect 2061 2548 2063 2551
rect 2087 2548 2089 2551
rect 2108 2548 2110 2551
rect 2128 2548 2130 2550
rect 2133 2548 2135 2551
rect 2151 2548 2153 2550
rect 2306 2555 2308 2559
rect 2334 2561 2336 2563
rect 2311 2555 2313 2558
rect 2201 2544 2203 2547
rect 2206 2545 2208 2547
rect 2202 2540 2203 2544
rect 2001 2526 2003 2540
rect 2017 2538 2019 2540
rect 2017 2526 2019 2528
rect 2033 2526 2035 2540
rect 2056 2535 2058 2540
rect 2061 2538 2063 2540
rect 2087 2538 2089 2540
rect 2052 2531 2058 2535
rect 2056 2526 2058 2531
rect 2061 2526 2063 2528
rect 2087 2526 2089 2528
rect 2108 2526 2110 2540
rect 2128 2535 2130 2540
rect 2133 2538 2135 2540
rect 2124 2531 2130 2535
rect 2128 2526 2130 2531
rect 2133 2526 2135 2528
rect 2151 2526 2153 2540
rect 2201 2535 2203 2540
rect 2206 2535 2208 2537
rect 2229 2531 2231 2553
rect 2280 2539 2282 2553
rect 2962 2555 2964 2558
rect 3006 2555 3008 2558
rect 3032 2555 3034 2558
rect 3078 2555 3080 2558
rect 3146 2555 3148 2559
rect 3174 2561 3176 2563
rect 3225 2561 3227 2563
rect 3151 2555 3153 2558
rect 2306 2544 2308 2547
rect 2311 2545 2313 2547
rect 2307 2540 2308 2544
rect 2306 2535 2308 2540
rect 2311 2535 2313 2537
rect 2280 2533 2282 2535
rect 2334 2531 2336 2553
rect 3032 2551 3033 2555
rect 2946 2548 2948 2550
rect 2962 2548 2964 2551
rect 2978 2548 2980 2550
rect 3001 2548 3003 2550
rect 3006 2548 3008 2551
rect 3032 2548 3034 2551
rect 3053 2548 3055 2551
rect 3073 2548 3075 2550
rect 3078 2548 3080 2551
rect 3096 2548 3098 2550
rect 3251 2555 3253 2559
rect 3279 2561 3281 2563
rect 3256 2555 3258 2558
rect 3146 2544 3148 2547
rect 3151 2545 3153 2547
rect 3147 2540 3148 2544
rect 2201 2529 2203 2531
rect 2206 2526 2208 2531
rect 2306 2529 2308 2531
rect 2229 2525 2231 2527
rect 2311 2526 2313 2531
rect 2334 2525 2336 2527
rect 2946 2526 2948 2540
rect 2962 2538 2964 2540
rect 2962 2526 2964 2528
rect 2978 2526 2980 2540
rect 3001 2535 3003 2540
rect 3006 2538 3008 2540
rect 3032 2538 3034 2540
rect 2997 2531 3003 2535
rect 3001 2526 3003 2531
rect 3006 2526 3008 2528
rect 3032 2526 3034 2528
rect 3053 2526 3055 2540
rect 3073 2535 3075 2540
rect 3078 2538 3080 2540
rect 3069 2531 3075 2535
rect 3073 2526 3075 2531
rect 3078 2526 3080 2528
rect 3096 2526 3098 2540
rect 3146 2535 3148 2540
rect 3151 2535 3153 2537
rect 3174 2531 3176 2553
rect 3225 2539 3227 2553
rect 3251 2544 3253 2547
rect 3256 2545 3258 2547
rect 3252 2540 3253 2544
rect 3251 2535 3253 2540
rect 3256 2535 3258 2537
rect 3225 2533 3227 2535
rect 3279 2531 3281 2553
rect 3146 2529 3148 2531
rect 3151 2526 3153 2531
rect 3251 2529 3253 2531
rect 3174 2525 3176 2527
rect 3256 2526 3258 2531
rect 3279 2525 3281 2527
rect 2001 2520 2003 2522
rect 2017 2518 2019 2522
rect 2033 2520 2035 2522
rect 2056 2520 2058 2522
rect 2018 2514 2019 2518
rect 2061 2517 2063 2522
rect 2087 2518 2089 2522
rect 2108 2520 2110 2522
rect 2128 2520 2130 2522
rect 2017 2511 2019 2514
rect 2062 2513 2063 2517
rect 2088 2514 2089 2518
rect 2133 2517 2135 2522
rect 2151 2520 2153 2522
rect 2946 2520 2948 2522
rect 2962 2518 2964 2522
rect 2978 2520 2980 2522
rect 3001 2520 3003 2522
rect 2061 2511 2063 2513
rect 2087 2510 2089 2514
rect 2134 2513 2135 2517
rect 2963 2514 2964 2518
rect 3006 2517 3008 2522
rect 3032 2518 3034 2522
rect 3053 2520 3055 2522
rect 3073 2520 3075 2522
rect 2133 2511 2135 2513
rect 2962 2511 2964 2514
rect 3007 2513 3008 2517
rect 3033 2514 3034 2518
rect 3078 2517 3080 2522
rect 3096 2520 3098 2522
rect 3006 2511 3008 2513
rect 3032 2510 3034 2514
rect 3079 2513 3080 2517
rect 3078 2511 3080 2513
rect 2017 2488 2019 2491
rect 2061 2489 2063 2491
rect 2018 2484 2019 2488
rect 2062 2485 2063 2489
rect 2087 2488 2089 2492
rect 2133 2489 2135 2491
rect 2001 2480 2003 2482
rect 2017 2480 2019 2484
rect 2033 2480 2035 2482
rect 2056 2480 2058 2482
rect 2061 2480 2063 2485
rect 2088 2484 2089 2488
rect 2134 2485 2135 2489
rect 2962 2488 2964 2491
rect 3006 2489 3008 2491
rect 2087 2480 2089 2484
rect 2108 2480 2110 2482
rect 2128 2480 2130 2482
rect 2133 2480 2135 2485
rect 2963 2484 2964 2488
rect 3007 2485 3008 2489
rect 3032 2488 3034 2492
rect 3078 2489 3080 2491
rect 2151 2480 2153 2482
rect 2201 2480 2203 2483
rect 2206 2480 2208 2483
rect 2306 2480 2308 2483
rect 2311 2480 2313 2483
rect 2946 2480 2948 2482
rect 2962 2480 2964 2484
rect 2978 2480 2980 2482
rect 3001 2480 3003 2482
rect 3006 2480 3008 2485
rect 3033 2484 3034 2488
rect 3079 2485 3080 2489
rect 3032 2480 3034 2484
rect 3053 2480 3055 2482
rect 3073 2480 3075 2482
rect 3078 2480 3080 2485
rect 3096 2480 3098 2482
rect 3146 2480 3148 2483
rect 3151 2480 3153 2483
rect 3251 2480 3253 2483
rect 3256 2480 3258 2483
rect 2001 2462 2003 2476
rect 2017 2474 2019 2476
rect 2017 2462 2019 2464
rect 2033 2462 2035 2476
rect 2056 2471 2058 2476
rect 2061 2474 2063 2476
rect 2087 2474 2089 2476
rect 2052 2467 2058 2471
rect 2056 2462 2058 2467
rect 2061 2462 2063 2464
rect 2087 2462 2089 2464
rect 2108 2462 2110 2476
rect 2128 2471 2130 2476
rect 2133 2474 2135 2476
rect 2124 2467 2130 2471
rect 2128 2462 2130 2467
rect 2133 2462 2135 2464
rect 2151 2462 2153 2476
rect 2201 2464 2203 2476
rect 2206 2474 2208 2476
rect 2206 2464 2208 2466
rect 2306 2464 2308 2476
rect 2311 2474 2313 2476
rect 2311 2464 2313 2466
rect 2946 2462 2948 2476
rect 2962 2474 2964 2476
rect 2962 2462 2964 2464
rect 2978 2462 2980 2476
rect 3001 2471 3003 2476
rect 3006 2474 3008 2476
rect 3032 2474 3034 2476
rect 2997 2467 3003 2471
rect 3001 2462 3003 2467
rect 3006 2462 3008 2464
rect 3032 2462 3034 2464
rect 3053 2462 3055 2476
rect 3073 2471 3075 2476
rect 3078 2474 3080 2476
rect 3069 2467 3075 2471
rect 3073 2462 3075 2467
rect 3078 2462 3080 2464
rect 3096 2462 3098 2476
rect 3146 2464 3148 2476
rect 3151 2474 3153 2476
rect 3151 2464 3153 2466
rect 3251 2464 3253 2476
rect 3256 2474 3258 2476
rect 3256 2464 3258 2466
rect 2201 2454 2203 2456
rect 2001 2452 2003 2454
rect 2017 2451 2019 2454
rect 2033 2452 2035 2454
rect 2056 2452 2058 2454
rect 2061 2451 2063 2454
rect 2087 2451 2089 2454
rect 2108 2451 2110 2454
rect 2128 2452 2130 2454
rect 2133 2451 2135 2454
rect 2151 2452 2153 2454
rect 2206 2451 2208 2456
rect 2306 2454 2308 2456
rect 2311 2451 2313 2456
rect 3146 2454 3148 2456
rect 2946 2452 2948 2454
rect 2087 2447 2088 2451
rect 2962 2451 2964 2454
rect 2978 2452 2980 2454
rect 3001 2452 3003 2454
rect 3006 2451 3008 2454
rect 3032 2451 3034 2454
rect 3053 2451 3055 2454
rect 3073 2452 3075 2454
rect 3078 2451 3080 2454
rect 3096 2452 3098 2454
rect 3151 2451 3153 2456
rect 3251 2454 3253 2456
rect 3256 2451 3258 2456
rect 3032 2447 3033 2451
rect 2017 2444 2019 2447
rect 2061 2444 2063 2447
rect 2087 2444 2089 2447
rect 2133 2444 2135 2447
rect 2962 2444 2964 2447
rect 3006 2444 3008 2447
rect 3032 2444 3034 2447
rect 3078 2444 3080 2447
rect 2017 2423 2019 2426
rect 2061 2423 2063 2426
rect 2087 2423 2089 2426
rect 2133 2423 2135 2426
rect 2201 2423 2203 2427
rect 2229 2429 2231 2431
rect 2256 2429 2258 2431
rect 2206 2423 2208 2426
rect 2087 2419 2088 2423
rect 2001 2416 2003 2418
rect 2017 2416 2019 2419
rect 2033 2416 2035 2418
rect 2056 2416 2058 2418
rect 2061 2416 2063 2419
rect 2087 2416 2089 2419
rect 2108 2416 2110 2419
rect 2128 2416 2130 2418
rect 2133 2416 2135 2419
rect 2151 2416 2153 2418
rect 2282 2423 2284 2427
rect 2310 2429 2312 2431
rect 2346 2429 2348 2431
rect 2287 2423 2289 2426
rect 2201 2412 2203 2415
rect 2206 2413 2208 2415
rect 2202 2408 2203 2412
rect 2001 2394 2003 2408
rect 2017 2406 2019 2408
rect 2017 2394 2019 2396
rect 2033 2394 2035 2408
rect 2056 2403 2058 2408
rect 2061 2406 2063 2408
rect 2087 2406 2089 2408
rect 2052 2399 2058 2403
rect 2056 2394 2058 2399
rect 2061 2394 2063 2396
rect 2087 2394 2089 2396
rect 2108 2394 2110 2408
rect 2128 2403 2130 2408
rect 2133 2406 2135 2408
rect 2124 2399 2130 2403
rect 2128 2394 2130 2399
rect 2133 2394 2135 2396
rect 2151 2394 2153 2408
rect 2201 2403 2203 2408
rect 2206 2403 2208 2405
rect 2229 2399 2231 2421
rect 2256 2407 2258 2421
rect 2372 2423 2374 2427
rect 2400 2429 2402 2431
rect 2377 2423 2379 2426
rect 2282 2412 2284 2415
rect 2287 2413 2289 2415
rect 2283 2408 2284 2412
rect 2282 2403 2284 2408
rect 2287 2403 2289 2405
rect 2256 2401 2258 2403
rect 2310 2399 2312 2421
rect 2346 2407 2348 2421
rect 2962 2423 2964 2426
rect 3006 2423 3008 2426
rect 3032 2423 3034 2426
rect 3078 2423 3080 2426
rect 3146 2423 3148 2427
rect 3174 2429 3176 2431
rect 3201 2429 3203 2431
rect 3151 2423 3153 2426
rect 2372 2412 2374 2415
rect 2377 2413 2379 2415
rect 2373 2408 2374 2412
rect 2372 2403 2374 2408
rect 2377 2403 2379 2405
rect 2346 2401 2348 2403
rect 2400 2399 2402 2421
rect 3032 2419 3033 2423
rect 2946 2416 2948 2418
rect 2962 2416 2964 2419
rect 2978 2416 2980 2418
rect 3001 2416 3003 2418
rect 3006 2416 3008 2419
rect 3032 2416 3034 2419
rect 3053 2416 3055 2419
rect 3073 2416 3075 2418
rect 3078 2416 3080 2419
rect 3096 2416 3098 2418
rect 3227 2423 3229 2427
rect 3255 2429 3257 2431
rect 3291 2429 3293 2431
rect 3232 2423 3234 2426
rect 3146 2412 3148 2415
rect 3151 2413 3153 2415
rect 3147 2408 3148 2412
rect 2201 2397 2203 2399
rect 2206 2394 2208 2399
rect 2282 2397 2284 2399
rect 2229 2393 2231 2395
rect 2287 2394 2289 2399
rect 2372 2397 2374 2399
rect 2310 2393 2312 2395
rect 2377 2394 2379 2399
rect 2400 2393 2402 2395
rect 2946 2394 2948 2408
rect 2962 2406 2964 2408
rect 2962 2394 2964 2396
rect 2978 2394 2980 2408
rect 3001 2403 3003 2408
rect 3006 2406 3008 2408
rect 3032 2406 3034 2408
rect 2997 2399 3003 2403
rect 3001 2394 3003 2399
rect 3006 2394 3008 2396
rect 3032 2394 3034 2396
rect 3053 2394 3055 2408
rect 3073 2403 3075 2408
rect 3078 2406 3080 2408
rect 3069 2399 3075 2403
rect 3073 2394 3075 2399
rect 3078 2394 3080 2396
rect 3096 2394 3098 2408
rect 3146 2403 3148 2408
rect 3151 2403 3153 2405
rect 3174 2399 3176 2421
rect 3201 2407 3203 2421
rect 3317 2423 3319 2427
rect 3345 2429 3347 2431
rect 3322 2423 3324 2426
rect 3227 2412 3229 2415
rect 3232 2413 3234 2415
rect 3228 2408 3229 2412
rect 3227 2403 3229 2408
rect 3232 2403 3234 2405
rect 3201 2401 3203 2403
rect 3255 2399 3257 2421
rect 3291 2407 3293 2421
rect 3317 2412 3319 2415
rect 3322 2413 3324 2415
rect 3318 2408 3319 2412
rect 3317 2403 3319 2408
rect 3322 2403 3324 2405
rect 3291 2401 3293 2403
rect 3345 2399 3347 2421
rect 3146 2397 3148 2399
rect 3151 2394 3153 2399
rect 3227 2397 3229 2399
rect 3174 2393 3176 2395
rect 3232 2394 3234 2399
rect 3317 2397 3319 2399
rect 3255 2393 3257 2395
rect 3322 2394 3324 2399
rect 3345 2393 3347 2395
rect 2001 2388 2003 2390
rect 2017 2386 2019 2390
rect 2033 2388 2035 2390
rect 2056 2388 2058 2390
rect 2018 2382 2019 2386
rect 2061 2385 2063 2390
rect 2087 2386 2089 2390
rect 2108 2388 2110 2390
rect 2128 2388 2130 2390
rect 2017 2379 2019 2382
rect 2062 2381 2063 2385
rect 2088 2382 2089 2386
rect 2133 2385 2135 2390
rect 2151 2388 2153 2390
rect 2946 2388 2948 2390
rect 2962 2386 2964 2390
rect 2978 2388 2980 2390
rect 3001 2388 3003 2390
rect 2061 2379 2063 2381
rect 2087 2378 2089 2382
rect 2134 2381 2135 2385
rect 2963 2382 2964 2386
rect 3006 2385 3008 2390
rect 3032 2386 3034 2390
rect 3053 2388 3055 2390
rect 3073 2388 3075 2390
rect 2133 2379 2135 2381
rect 2962 2379 2964 2382
rect 3007 2381 3008 2385
rect 3033 2382 3034 2386
rect 3078 2385 3080 2390
rect 3096 2388 3098 2390
rect 3006 2379 3008 2381
rect 3032 2378 3034 2382
rect 3079 2381 3080 2385
rect 3078 2379 3080 2381
rect 2017 2356 2019 2359
rect 2061 2357 2063 2359
rect 2018 2352 2019 2356
rect 2062 2353 2063 2357
rect 2087 2356 2089 2360
rect 2133 2357 2135 2359
rect 2001 2348 2003 2350
rect 2017 2348 2019 2352
rect 2033 2348 2035 2350
rect 2056 2348 2058 2350
rect 2061 2348 2063 2353
rect 2088 2352 2089 2356
rect 2134 2353 2135 2357
rect 2962 2356 2964 2359
rect 3006 2357 3008 2359
rect 2087 2348 2089 2352
rect 2108 2348 2110 2350
rect 2128 2348 2130 2350
rect 2133 2348 2135 2353
rect 2963 2352 2964 2356
rect 3007 2353 3008 2357
rect 3032 2356 3034 2360
rect 3078 2357 3080 2359
rect 2151 2348 2153 2350
rect 2946 2348 2948 2350
rect 2962 2348 2964 2352
rect 2978 2348 2980 2350
rect 3001 2348 3003 2350
rect 3006 2348 3008 2353
rect 3033 2352 3034 2356
rect 3079 2353 3080 2357
rect 3032 2348 3034 2352
rect 3053 2348 3055 2350
rect 3073 2348 3075 2350
rect 3078 2348 3080 2353
rect 3096 2348 3098 2350
rect 2201 2345 2203 2348
rect 2206 2345 2208 2348
rect 2282 2345 2284 2348
rect 2287 2345 2289 2348
rect 2372 2345 2374 2348
rect 2377 2345 2379 2348
rect 2001 2330 2003 2344
rect 2017 2342 2019 2344
rect 2017 2330 2019 2332
rect 2033 2330 2035 2344
rect 2056 2339 2058 2344
rect 2061 2342 2063 2344
rect 2087 2342 2089 2344
rect 2052 2335 2058 2339
rect 2056 2330 2058 2335
rect 2061 2330 2063 2332
rect 2087 2330 2089 2332
rect 2108 2330 2110 2344
rect 2128 2339 2130 2344
rect 2133 2342 2135 2344
rect 2124 2335 2130 2339
rect 2128 2330 2130 2335
rect 2133 2330 2135 2332
rect 2151 2330 2153 2344
rect 3146 2345 3148 2348
rect 3151 2345 3153 2348
rect 3227 2345 3229 2348
rect 3232 2345 3234 2348
rect 3317 2345 3319 2348
rect 3322 2345 3324 2348
rect 2201 2329 2203 2341
rect 2206 2339 2208 2341
rect 2206 2329 2208 2331
rect 2282 2329 2284 2341
rect 2287 2339 2289 2341
rect 2287 2329 2289 2331
rect 2372 2329 2374 2341
rect 2377 2339 2379 2341
rect 2377 2329 2379 2331
rect 2946 2330 2948 2344
rect 2962 2342 2964 2344
rect 2962 2330 2964 2332
rect 2978 2330 2980 2344
rect 3001 2339 3003 2344
rect 3006 2342 3008 2344
rect 3032 2342 3034 2344
rect 2997 2335 3003 2339
rect 3001 2330 3003 2335
rect 3006 2330 3008 2332
rect 3032 2330 3034 2332
rect 3053 2330 3055 2344
rect 3073 2339 3075 2344
rect 3078 2342 3080 2344
rect 3069 2335 3075 2339
rect 3073 2330 3075 2335
rect 3078 2330 3080 2332
rect 3096 2330 3098 2344
rect 2001 2320 2003 2322
rect 2017 2319 2019 2322
rect 2033 2320 2035 2322
rect 2056 2320 2058 2322
rect 2061 2319 2063 2322
rect 2087 2319 2089 2322
rect 2108 2319 2110 2322
rect 2128 2320 2130 2322
rect 2133 2319 2135 2322
rect 2151 2320 2153 2322
rect 3146 2329 3148 2341
rect 3151 2339 3153 2341
rect 3151 2329 3153 2331
rect 3227 2329 3229 2341
rect 3232 2339 3234 2341
rect 3232 2329 3234 2331
rect 3317 2329 3319 2341
rect 3322 2339 3324 2341
rect 3322 2329 3324 2331
rect 2201 2319 2203 2321
rect 2087 2315 2088 2319
rect 2206 2316 2208 2321
rect 2282 2319 2284 2321
rect 2287 2316 2289 2321
rect 2372 2319 2374 2321
rect 2377 2316 2379 2321
rect 2946 2320 2948 2322
rect 2017 2312 2019 2315
rect 2061 2312 2063 2315
rect 2087 2312 2089 2315
rect 2133 2312 2135 2315
rect 2962 2319 2964 2322
rect 2978 2320 2980 2322
rect 3001 2320 3003 2322
rect 3006 2319 3008 2322
rect 3032 2319 3034 2322
rect 3053 2319 3055 2322
rect 3073 2320 3075 2322
rect 3078 2319 3080 2322
rect 3096 2320 3098 2322
rect 3146 2319 3148 2321
rect 3032 2315 3033 2319
rect 3151 2316 3153 2321
rect 3227 2319 3229 2321
rect 3232 2316 3234 2321
rect 3317 2319 3319 2321
rect 3322 2316 3324 2321
rect 2962 2312 2964 2315
rect 3006 2312 3008 2315
rect 3032 2312 3034 2315
rect 3078 2312 3080 2315
rect 2017 2291 2019 2294
rect 2061 2291 2063 2294
rect 2087 2291 2089 2294
rect 2133 2291 2135 2294
rect 2201 2291 2203 2295
rect 2229 2297 2231 2299
rect 2206 2291 2208 2294
rect 2087 2287 2088 2291
rect 2001 2284 2003 2286
rect 2017 2284 2019 2287
rect 2033 2284 2035 2286
rect 2056 2284 2058 2286
rect 2061 2284 2063 2287
rect 2087 2284 2089 2287
rect 2108 2284 2110 2287
rect 2128 2284 2130 2286
rect 2133 2284 2135 2287
rect 2151 2284 2153 2286
rect 2962 2291 2964 2294
rect 3006 2291 3008 2294
rect 3032 2291 3034 2294
rect 3078 2291 3080 2294
rect 3146 2291 3148 2295
rect 3174 2297 3176 2299
rect 3151 2291 3153 2294
rect 2201 2280 2203 2283
rect 2206 2281 2208 2283
rect 2202 2276 2203 2280
rect 2001 2262 2003 2276
rect 2017 2274 2019 2276
rect 2017 2262 2019 2264
rect 2033 2262 2035 2276
rect 2056 2271 2058 2276
rect 2061 2274 2063 2276
rect 2087 2274 2089 2276
rect 2052 2267 2058 2271
rect 2056 2262 2058 2267
rect 2061 2262 2063 2264
rect 2087 2262 2089 2264
rect 2108 2262 2110 2276
rect 2128 2271 2130 2276
rect 2133 2274 2135 2276
rect 2124 2267 2130 2271
rect 2128 2262 2130 2267
rect 2133 2262 2135 2264
rect 2151 2262 2153 2276
rect 2201 2271 2203 2276
rect 2206 2271 2208 2273
rect 2229 2267 2231 2289
rect 3032 2287 3033 2291
rect 2946 2284 2948 2286
rect 2962 2284 2964 2287
rect 2978 2284 2980 2286
rect 3001 2284 3003 2286
rect 3006 2284 3008 2287
rect 3032 2284 3034 2287
rect 3053 2284 3055 2287
rect 3073 2284 3075 2286
rect 3078 2284 3080 2287
rect 3096 2284 3098 2286
rect 3146 2280 3148 2283
rect 3151 2281 3153 2283
rect 3147 2276 3148 2280
rect 2201 2265 2203 2267
rect 2206 2262 2208 2267
rect 2229 2261 2231 2263
rect 2946 2262 2948 2276
rect 2962 2274 2964 2276
rect 2962 2262 2964 2264
rect 2978 2262 2980 2276
rect 3001 2271 3003 2276
rect 3006 2274 3008 2276
rect 3032 2274 3034 2276
rect 2997 2267 3003 2271
rect 3001 2262 3003 2267
rect 3006 2262 3008 2264
rect 3032 2262 3034 2264
rect 3053 2262 3055 2276
rect 3073 2271 3075 2276
rect 3078 2274 3080 2276
rect 3069 2267 3075 2271
rect 3073 2262 3075 2267
rect 3078 2262 3080 2264
rect 3096 2262 3098 2276
rect 3146 2271 3148 2276
rect 3151 2271 3153 2273
rect 3174 2267 3176 2289
rect 3146 2265 3148 2267
rect 3151 2262 3153 2267
rect 3174 2261 3176 2263
rect 2001 2256 2003 2258
rect 2017 2254 2019 2258
rect 2033 2256 2035 2258
rect 2056 2256 2058 2258
rect 2018 2250 2019 2254
rect 2061 2253 2063 2258
rect 2087 2254 2089 2258
rect 2108 2256 2110 2258
rect 2128 2256 2130 2258
rect 2017 2247 2019 2250
rect 2062 2249 2063 2253
rect 2088 2250 2089 2254
rect 2133 2253 2135 2258
rect 2151 2256 2153 2258
rect 2946 2256 2948 2258
rect 2962 2254 2964 2258
rect 2978 2256 2980 2258
rect 3001 2256 3003 2258
rect 2061 2247 2063 2249
rect 2087 2246 2089 2250
rect 2134 2249 2135 2253
rect 2963 2250 2964 2254
rect 3006 2253 3008 2258
rect 3032 2254 3034 2258
rect 3053 2256 3055 2258
rect 3073 2256 3075 2258
rect 2133 2247 2135 2249
rect 2962 2247 2964 2250
rect 3007 2249 3008 2253
rect 3033 2250 3034 2254
rect 3078 2253 3080 2258
rect 3096 2256 3098 2258
rect 3006 2247 3008 2249
rect 3032 2246 3034 2250
rect 3079 2249 3080 2253
rect 3078 2247 3080 2249
rect 1512 2229 1514 2231
rect 1517 2229 1519 2232
rect 1533 2229 1535 2231
rect 1549 2229 1551 2231
rect 1554 2229 1556 2232
rect 1575 2229 1577 2232
rect 1591 2229 1593 2232
rect 1607 2229 1609 2231
rect 1612 2229 1614 2232
rect 1628 2229 1630 2231
rect 1644 2229 1646 2231
rect 1649 2229 1651 2232
rect 1665 2229 1667 2231
rect 1681 2229 1683 2231
rect 1686 2229 1688 2232
rect 1707 2229 1709 2232
rect 1723 2229 1725 2232
rect 1739 2229 1741 2231
rect 1744 2229 1746 2232
rect 1760 2229 1762 2231
rect 1776 2229 1778 2231
rect 1781 2229 1783 2232
rect 1797 2229 1799 2231
rect 1813 2229 1815 2231
rect 1818 2229 1820 2232
rect 1839 2229 1841 2232
rect 1855 2229 1857 2232
rect 1871 2229 1873 2231
rect 1876 2229 1878 2232
rect 1892 2229 1894 2231
rect 2457 2229 2459 2231
rect 2462 2229 2464 2232
rect 2478 2229 2480 2231
rect 2494 2229 2496 2231
rect 2499 2229 2501 2232
rect 2520 2229 2522 2232
rect 2536 2229 2538 2232
rect 2552 2229 2554 2231
rect 2557 2229 2559 2232
rect 2573 2229 2575 2231
rect 2589 2229 2591 2231
rect 2594 2229 2596 2232
rect 2610 2229 2612 2231
rect 2626 2229 2628 2231
rect 2631 2229 2633 2232
rect 2652 2229 2654 2232
rect 2668 2229 2670 2232
rect 2684 2229 2686 2231
rect 2689 2229 2691 2232
rect 2705 2229 2707 2231
rect 2721 2229 2723 2231
rect 2726 2229 2728 2232
rect 2742 2229 2744 2231
rect 2758 2229 2760 2231
rect 2763 2229 2765 2232
rect 2784 2229 2786 2232
rect 2800 2229 2802 2232
rect 2816 2229 2818 2231
rect 2821 2229 2823 2232
rect 2837 2229 2839 2231
rect 2017 2224 2019 2227
rect 2061 2225 2063 2227
rect 1512 2216 1514 2221
rect 1517 2219 1519 2221
rect 1512 2202 1514 2212
rect 1517 2202 1519 2209
rect 1533 2202 1535 2221
rect 1549 2212 1551 2221
rect 1554 2219 1556 2221
rect 1575 2219 1577 2221
rect 1591 2218 1593 2221
rect 1549 2202 1551 2205
rect 1554 2202 1556 2204
rect 1575 2202 1577 2204
rect 1591 2202 1593 2214
rect 1607 2212 1609 2221
rect 1612 2219 1614 2221
rect 1607 2202 1609 2205
rect 1612 2202 1614 2204
rect 1628 2202 1630 2221
rect 1644 2218 1646 2221
rect 1649 2219 1651 2221
rect 1644 2202 1646 2214
rect 1649 2202 1651 2209
rect 1665 2202 1667 2221
rect 1681 2212 1683 2221
rect 1686 2219 1688 2221
rect 1707 2219 1709 2221
rect 1723 2218 1725 2221
rect 1681 2202 1683 2205
rect 1686 2202 1688 2204
rect 1707 2202 1709 2204
rect 1723 2202 1725 2214
rect 1739 2212 1741 2221
rect 1744 2219 1746 2221
rect 1739 2202 1741 2205
rect 1744 2202 1746 2204
rect 1760 2202 1762 2221
rect 1776 2218 1778 2221
rect 1781 2219 1783 2221
rect 1776 2202 1778 2214
rect 1781 2202 1783 2209
rect 1797 2202 1799 2221
rect 1813 2212 1815 2221
rect 1818 2219 1820 2221
rect 1839 2219 1841 2221
rect 1855 2218 1857 2221
rect 1813 2202 1815 2205
rect 1818 2202 1820 2204
rect 1839 2202 1841 2204
rect 1855 2202 1857 2214
rect 1871 2212 1873 2221
rect 1876 2219 1878 2221
rect 1892 2213 1894 2221
rect 2018 2220 2019 2224
rect 2062 2221 2063 2225
rect 2087 2224 2089 2228
rect 2133 2225 2135 2227
rect 2001 2216 2003 2218
rect 2017 2216 2019 2220
rect 2033 2216 2035 2218
rect 2056 2216 2058 2218
rect 2061 2216 2063 2221
rect 2088 2220 2089 2224
rect 2134 2221 2135 2225
rect 2278 2224 2280 2227
rect 2322 2225 2324 2227
rect 2087 2216 2089 2220
rect 2108 2216 2110 2218
rect 2128 2216 2130 2218
rect 2133 2216 2135 2221
rect 2279 2220 2280 2224
rect 2323 2221 2324 2225
rect 2348 2224 2350 2228
rect 2394 2225 2396 2227
rect 2151 2216 2153 2218
rect 2235 2216 2237 2219
rect 2253 2216 2255 2219
rect 2278 2216 2280 2220
rect 2294 2216 2296 2218
rect 2317 2216 2319 2218
rect 2322 2216 2324 2221
rect 2349 2220 2350 2224
rect 2395 2221 2396 2225
rect 2962 2224 2964 2227
rect 3006 2225 3008 2227
rect 2348 2216 2350 2220
rect 2369 2216 2371 2218
rect 2389 2216 2391 2218
rect 2394 2216 2396 2221
rect 2412 2216 2414 2218
rect 2457 2216 2459 2221
rect 2462 2219 2464 2221
rect 1871 2202 1873 2205
rect 1876 2202 1878 2204
rect 1892 2202 1894 2209
rect 2001 2198 2003 2212
rect 2017 2210 2019 2212
rect 2017 2198 2019 2200
rect 2033 2198 2035 2212
rect 2056 2207 2058 2212
rect 2061 2210 2063 2212
rect 2087 2210 2089 2212
rect 2052 2203 2058 2207
rect 2056 2198 2058 2203
rect 2061 2198 2063 2200
rect 2087 2198 2089 2200
rect 2108 2198 2110 2212
rect 2128 2207 2130 2212
rect 2133 2210 2135 2212
rect 2124 2203 2130 2207
rect 2128 2198 2130 2203
rect 2133 2198 2135 2200
rect 2151 2198 2153 2212
rect 2201 2209 2203 2212
rect 2206 2209 2208 2212
rect 2235 2207 2237 2212
rect 1512 2196 1514 2198
rect 1517 2195 1519 2198
rect 1533 2196 1535 2198
rect 1549 2196 1551 2198
rect 1554 2193 1556 2198
rect 1575 2193 1577 2198
rect 1591 2196 1593 2198
rect 1607 2196 1609 2198
rect 1612 2193 1614 2198
rect 1628 2196 1630 2198
rect 1644 2196 1646 2198
rect 1649 2195 1651 2198
rect 1665 2196 1667 2198
rect 1681 2196 1683 2198
rect 1686 2193 1688 2198
rect 1707 2193 1709 2198
rect 1723 2196 1725 2198
rect 1739 2196 1741 2198
rect 1744 2193 1746 2198
rect 1760 2196 1762 2198
rect 1776 2196 1778 2198
rect 1781 2195 1783 2198
rect 1797 2196 1799 2198
rect 1813 2196 1815 2198
rect 1818 2193 1820 2198
rect 1839 2193 1841 2198
rect 1855 2196 1857 2198
rect 1871 2196 1873 2198
rect 1876 2193 1878 2198
rect 1892 2196 1894 2198
rect 2201 2193 2203 2205
rect 2206 2203 2208 2205
rect 2235 2198 2237 2203
rect 2253 2198 2255 2212
rect 2278 2210 2280 2212
rect 2278 2198 2280 2200
rect 2294 2198 2296 2212
rect 2317 2207 2319 2212
rect 2322 2210 2324 2212
rect 2348 2210 2350 2212
rect 2313 2203 2319 2207
rect 2317 2198 2319 2203
rect 2322 2198 2324 2200
rect 2348 2198 2350 2200
rect 2369 2198 2371 2212
rect 2389 2207 2391 2212
rect 2394 2210 2396 2212
rect 2385 2203 2391 2207
rect 2389 2198 2391 2203
rect 2394 2198 2396 2200
rect 2412 2198 2414 2212
rect 2457 2202 2459 2212
rect 2462 2202 2464 2209
rect 2478 2202 2480 2221
rect 2494 2212 2496 2221
rect 2499 2219 2501 2221
rect 2520 2219 2522 2221
rect 2536 2218 2538 2221
rect 2494 2202 2496 2205
rect 2499 2202 2501 2204
rect 2520 2202 2522 2204
rect 2536 2202 2538 2214
rect 2552 2212 2554 2221
rect 2557 2219 2559 2221
rect 2552 2202 2554 2205
rect 2557 2202 2559 2204
rect 2573 2202 2575 2221
rect 2589 2218 2591 2221
rect 2594 2219 2596 2221
rect 2589 2202 2591 2214
rect 2594 2202 2596 2209
rect 2610 2202 2612 2221
rect 2626 2212 2628 2221
rect 2631 2219 2633 2221
rect 2652 2219 2654 2221
rect 2668 2218 2670 2221
rect 2626 2202 2628 2205
rect 2631 2202 2633 2204
rect 2652 2202 2654 2204
rect 2668 2202 2670 2214
rect 2684 2212 2686 2221
rect 2689 2219 2691 2221
rect 2684 2202 2686 2205
rect 2689 2202 2691 2204
rect 2705 2202 2707 2221
rect 2721 2218 2723 2221
rect 2726 2219 2728 2221
rect 2721 2202 2723 2214
rect 2726 2202 2728 2209
rect 2742 2202 2744 2221
rect 2758 2212 2760 2221
rect 2763 2219 2765 2221
rect 2784 2219 2786 2221
rect 2800 2218 2802 2221
rect 2758 2202 2760 2205
rect 2763 2202 2765 2204
rect 2784 2202 2786 2204
rect 2800 2202 2802 2214
rect 2816 2212 2818 2221
rect 2821 2219 2823 2221
rect 2837 2213 2839 2221
rect 2963 2220 2964 2224
rect 3007 2221 3008 2225
rect 3032 2224 3034 2228
rect 3078 2225 3080 2227
rect 2946 2216 2948 2218
rect 2962 2216 2964 2220
rect 2978 2216 2980 2218
rect 3001 2216 3003 2218
rect 3006 2216 3008 2221
rect 3033 2220 3034 2224
rect 3079 2221 3080 2225
rect 3223 2224 3225 2227
rect 3267 2225 3269 2227
rect 3032 2216 3034 2220
rect 3053 2216 3055 2218
rect 3073 2216 3075 2218
rect 3078 2216 3080 2221
rect 3224 2220 3225 2224
rect 3268 2221 3269 2225
rect 3293 2224 3295 2228
rect 3339 2225 3341 2227
rect 3096 2216 3098 2218
rect 3180 2216 3182 2219
rect 3198 2216 3200 2219
rect 3223 2216 3225 2220
rect 3239 2216 3241 2218
rect 3262 2216 3264 2218
rect 3267 2216 3269 2221
rect 3294 2220 3295 2224
rect 3340 2221 3341 2225
rect 3293 2216 3295 2220
rect 3314 2216 3316 2218
rect 3334 2216 3336 2218
rect 3339 2216 3341 2221
rect 3357 2216 3359 2218
rect 2816 2202 2818 2205
rect 2821 2202 2823 2204
rect 2837 2202 2839 2209
rect 2946 2198 2948 2212
rect 2962 2210 2964 2212
rect 2962 2198 2964 2200
rect 2978 2198 2980 2212
rect 3001 2207 3003 2212
rect 3006 2210 3008 2212
rect 3032 2210 3034 2212
rect 2997 2203 3003 2207
rect 3001 2198 3003 2203
rect 3006 2198 3008 2200
rect 3032 2198 3034 2200
rect 3053 2198 3055 2212
rect 3073 2207 3075 2212
rect 3078 2210 3080 2212
rect 3069 2203 3075 2207
rect 3073 2198 3075 2203
rect 3078 2198 3080 2200
rect 3096 2198 3098 2212
rect 3146 2209 3148 2212
rect 3151 2209 3153 2212
rect 3180 2207 3182 2212
rect 2206 2193 2208 2195
rect 2001 2188 2003 2190
rect 2017 2187 2019 2190
rect 2033 2188 2035 2190
rect 2056 2188 2058 2190
rect 2061 2187 2063 2190
rect 2087 2187 2089 2190
rect 2108 2187 2110 2190
rect 2128 2188 2130 2190
rect 2133 2187 2135 2190
rect 2151 2188 2153 2190
rect 2087 2183 2088 2187
rect 2457 2196 2459 2198
rect 2462 2195 2464 2198
rect 2478 2196 2480 2198
rect 2494 2196 2496 2198
rect 2499 2193 2501 2198
rect 2520 2193 2522 2198
rect 2536 2196 2538 2198
rect 2552 2196 2554 2198
rect 2557 2193 2559 2198
rect 2573 2196 2575 2198
rect 2589 2196 2591 2198
rect 2235 2187 2237 2190
rect 2201 2183 2203 2185
rect 2017 2180 2019 2183
rect 2061 2180 2063 2183
rect 2087 2180 2089 2183
rect 2133 2180 2135 2183
rect 2206 2180 2208 2185
rect 1627 2158 1629 2161
rect 1651 2158 1653 2161
rect 1627 2152 1629 2154
rect 1651 2152 1653 2154
rect 2253 2148 2255 2190
rect 2278 2187 2280 2190
rect 2294 2188 2296 2190
rect 2317 2188 2319 2190
rect 2322 2187 2324 2190
rect 2348 2187 2350 2190
rect 2369 2187 2371 2190
rect 2389 2188 2391 2190
rect 2394 2187 2396 2190
rect 2412 2188 2414 2190
rect 2594 2195 2596 2198
rect 2610 2196 2612 2198
rect 2626 2196 2628 2198
rect 2631 2193 2633 2198
rect 2652 2193 2654 2198
rect 2668 2196 2670 2198
rect 2684 2196 2686 2198
rect 2689 2193 2691 2198
rect 2705 2196 2707 2198
rect 2721 2196 2723 2198
rect 2726 2195 2728 2198
rect 2742 2196 2744 2198
rect 2758 2196 2760 2198
rect 2763 2193 2765 2198
rect 2784 2193 2786 2198
rect 2800 2196 2802 2198
rect 2816 2196 2818 2198
rect 2821 2193 2823 2198
rect 2837 2196 2839 2198
rect 3146 2193 3148 2205
rect 3151 2203 3153 2205
rect 3180 2198 3182 2203
rect 3198 2198 3200 2212
rect 3223 2210 3225 2212
rect 3223 2198 3225 2200
rect 3239 2198 3241 2212
rect 3262 2207 3264 2212
rect 3267 2210 3269 2212
rect 3293 2210 3295 2212
rect 3258 2203 3264 2207
rect 3262 2198 3264 2203
rect 3267 2198 3269 2200
rect 3293 2198 3295 2200
rect 3314 2198 3316 2212
rect 3334 2207 3336 2212
rect 3339 2210 3341 2212
rect 3330 2203 3336 2207
rect 3334 2198 3336 2203
rect 3339 2198 3341 2200
rect 3357 2198 3359 2212
rect 3151 2193 3153 2195
rect 2946 2188 2948 2190
rect 2962 2187 2964 2190
rect 2978 2188 2980 2190
rect 3001 2188 3003 2190
rect 3006 2187 3008 2190
rect 3032 2187 3034 2190
rect 3053 2187 3055 2190
rect 3073 2188 3075 2190
rect 3078 2187 3080 2190
rect 3096 2188 3098 2190
rect 2348 2183 2349 2187
rect 2278 2180 2280 2183
rect 2322 2180 2324 2183
rect 2348 2180 2350 2183
rect 2394 2180 2396 2183
rect 3032 2183 3033 2187
rect 3180 2187 3182 2190
rect 3146 2183 3148 2185
rect 2962 2180 2964 2183
rect 3006 2180 3008 2183
rect 3032 2180 3034 2183
rect 3078 2180 3080 2183
rect 3151 2180 3153 2185
rect 2572 2158 2574 2161
rect 2596 2158 2598 2161
rect 2421 2156 2424 2158
rect 2428 2156 2431 2158
rect 2572 2152 2574 2154
rect 2596 2152 2598 2154
rect 3198 2152 3200 2190
rect 3223 2187 3225 2190
rect 3239 2188 3241 2190
rect 3262 2188 3264 2190
rect 3267 2187 3269 2190
rect 3293 2187 3295 2190
rect 3314 2187 3316 2190
rect 3334 2188 3336 2190
rect 3339 2187 3341 2190
rect 3357 2188 3359 2190
rect 3293 2183 3294 2187
rect 3223 2180 3225 2183
rect 3267 2180 3269 2183
rect 3293 2180 3295 2183
rect 3339 2180 3341 2183
rect 3366 2156 3369 2158
rect 3373 2156 3376 2158
rect 1647 2145 1649 2147
rect 2592 2145 2594 2147
rect 1647 2138 1649 2141
rect 2592 2138 2594 2141
rect 1636 2127 1638 2129
rect 1642 2127 1661 2129
rect 2581 2127 2583 2129
rect 2587 2127 2606 2129
rect 1627 2122 1629 2124
rect 1651 2122 1653 2124
rect 2572 2122 2574 2124
rect 2596 2122 2598 2124
rect 1627 2115 1629 2118
rect 1651 2115 1653 2118
rect 2295 2117 2297 2119
rect 2300 2117 2302 2120
rect 2316 2117 2318 2119
rect 2332 2117 2334 2119
rect 2337 2117 2339 2120
rect 2358 2117 2360 2120
rect 2374 2117 2376 2120
rect 2390 2117 2392 2119
rect 2395 2117 2397 2120
rect 2411 2117 2413 2119
rect 2572 2115 2574 2118
rect 2596 2115 2598 2118
rect 3240 2117 3242 2119
rect 3245 2117 3247 2120
rect 3261 2117 3263 2119
rect 3277 2117 3279 2119
rect 3282 2117 3284 2120
rect 3303 2117 3305 2120
rect 3319 2117 3321 2120
rect 3335 2117 3337 2119
rect 3340 2117 3342 2120
rect 3356 2117 3358 2119
rect 2295 2104 2297 2109
rect 2300 2107 2302 2109
rect 2295 2090 2297 2100
rect 2300 2090 2302 2097
rect 2316 2090 2318 2109
rect 2332 2100 2334 2109
rect 2337 2107 2339 2109
rect 2358 2107 2360 2109
rect 2374 2106 2376 2109
rect 2332 2090 2334 2093
rect 2337 2090 2339 2092
rect 2358 2090 2360 2092
rect 2374 2090 2376 2102
rect 2390 2100 2392 2109
rect 2395 2107 2397 2109
rect 2390 2090 2392 2093
rect 2395 2090 2397 2092
rect 2411 2090 2413 2109
rect 3240 2104 3242 2109
rect 3245 2107 3247 2109
rect 3240 2090 3242 2100
rect 3245 2090 3247 2097
rect 3261 2090 3263 2109
rect 3277 2100 3279 2109
rect 3282 2107 3284 2109
rect 3303 2107 3305 2109
rect 3319 2106 3321 2109
rect 3277 2090 3279 2093
rect 3282 2090 3284 2092
rect 3303 2090 3305 2092
rect 3319 2090 3321 2102
rect 3335 2100 3337 2109
rect 3340 2107 3342 2109
rect 3335 2090 3337 2093
rect 3340 2090 3342 2092
rect 3356 2090 3358 2109
rect 1512 2087 1514 2089
rect 1517 2087 1519 2090
rect 1533 2087 1535 2089
rect 1549 2087 1551 2089
rect 1554 2087 1556 2090
rect 1575 2087 1577 2090
rect 1591 2087 1593 2090
rect 1607 2087 1609 2089
rect 1612 2087 1614 2090
rect 1628 2087 1630 2089
rect 1644 2087 1646 2089
rect 1649 2087 1651 2090
rect 1665 2087 1667 2089
rect 1681 2087 1683 2089
rect 1686 2087 1688 2090
rect 1707 2087 1709 2090
rect 1723 2087 1725 2090
rect 1739 2087 1741 2089
rect 1744 2087 1746 2090
rect 1760 2087 1762 2089
rect 1776 2087 1778 2089
rect 1781 2087 1783 2090
rect 1797 2087 1799 2089
rect 1813 2087 1815 2089
rect 1818 2087 1820 2090
rect 1839 2087 1841 2090
rect 1855 2087 1857 2090
rect 1871 2087 1873 2089
rect 1876 2087 1878 2090
rect 1892 2087 1894 2089
rect 2457 2087 2459 2089
rect 2462 2087 2464 2090
rect 2478 2087 2480 2089
rect 2494 2087 2496 2089
rect 2499 2087 2501 2090
rect 2520 2087 2522 2090
rect 2536 2087 2538 2090
rect 2552 2087 2554 2089
rect 2557 2087 2559 2090
rect 2573 2087 2575 2089
rect 2589 2087 2591 2089
rect 2594 2087 2596 2090
rect 2610 2087 2612 2089
rect 2626 2087 2628 2089
rect 2631 2087 2633 2090
rect 2652 2087 2654 2090
rect 2668 2087 2670 2090
rect 2684 2087 2686 2089
rect 2689 2087 2691 2090
rect 2705 2087 2707 2089
rect 2721 2087 2723 2089
rect 2726 2087 2728 2090
rect 2742 2087 2744 2089
rect 2758 2087 2760 2089
rect 2763 2087 2765 2090
rect 2784 2087 2786 2090
rect 2800 2087 2802 2090
rect 2816 2087 2818 2089
rect 2821 2087 2823 2090
rect 2837 2087 2839 2089
rect 2295 2084 2297 2086
rect 2300 2083 2302 2086
rect 2316 2084 2318 2086
rect 2332 2084 2334 2086
rect 2337 2081 2339 2086
rect 2358 2081 2360 2086
rect 2374 2084 2376 2086
rect 2390 2084 2392 2086
rect 2395 2081 2397 2086
rect 2411 2084 2413 2086
rect 1512 2074 1514 2079
rect 1517 2077 1519 2079
rect 1512 2060 1514 2070
rect 1517 2060 1519 2067
rect 1533 2060 1535 2079
rect 1549 2070 1551 2079
rect 1554 2077 1556 2079
rect 1575 2077 1577 2079
rect 1591 2076 1593 2079
rect 1549 2060 1551 2063
rect 1554 2060 1556 2062
rect 1575 2060 1577 2062
rect 1591 2060 1593 2072
rect 1607 2070 1609 2079
rect 1612 2077 1614 2079
rect 1607 2060 1609 2063
rect 1612 2060 1614 2062
rect 1628 2060 1630 2079
rect 1644 2076 1646 2079
rect 1649 2077 1651 2079
rect 1644 2060 1646 2072
rect 1649 2060 1651 2067
rect 1665 2060 1667 2079
rect 1681 2070 1683 2079
rect 1686 2077 1688 2079
rect 1707 2077 1709 2079
rect 1723 2076 1725 2079
rect 1681 2060 1683 2063
rect 1686 2060 1688 2062
rect 1707 2060 1709 2062
rect 1723 2060 1725 2072
rect 1739 2070 1741 2079
rect 1744 2077 1746 2079
rect 1739 2060 1741 2063
rect 1744 2060 1746 2062
rect 1760 2060 1762 2079
rect 1776 2076 1778 2079
rect 1781 2077 1783 2079
rect 1776 2060 1778 2072
rect 1781 2060 1783 2067
rect 1797 2060 1799 2079
rect 1813 2070 1815 2079
rect 1818 2077 1820 2079
rect 1839 2077 1841 2079
rect 1855 2076 1857 2079
rect 1813 2060 1815 2063
rect 1818 2060 1820 2062
rect 1839 2060 1841 2062
rect 1855 2060 1857 2072
rect 1871 2070 1873 2079
rect 1876 2077 1878 2079
rect 1892 2071 1894 2079
rect 3240 2084 3242 2086
rect 3245 2083 3247 2086
rect 3261 2084 3263 2086
rect 3277 2084 3279 2086
rect 3282 2081 3284 2086
rect 3303 2081 3305 2086
rect 3319 2084 3321 2086
rect 3335 2084 3337 2086
rect 3340 2081 3342 2086
rect 3356 2084 3358 2086
rect 2457 2074 2459 2079
rect 2462 2077 2464 2079
rect 1871 2060 1873 2063
rect 1876 2060 1878 2062
rect 1892 2060 1894 2067
rect 2457 2060 2459 2070
rect 2462 2060 2464 2067
rect 2478 2060 2480 2079
rect 2494 2070 2496 2079
rect 2499 2077 2501 2079
rect 2520 2077 2522 2079
rect 2536 2076 2538 2079
rect 2494 2060 2496 2063
rect 2499 2060 2501 2062
rect 2520 2060 2522 2062
rect 2536 2060 2538 2072
rect 2552 2070 2554 2079
rect 2557 2077 2559 2079
rect 2552 2060 2554 2063
rect 2557 2060 2559 2062
rect 2573 2060 2575 2079
rect 2589 2076 2591 2079
rect 2594 2077 2596 2079
rect 2589 2060 2591 2072
rect 2594 2060 2596 2067
rect 2610 2060 2612 2079
rect 2626 2070 2628 2079
rect 2631 2077 2633 2079
rect 2652 2077 2654 2079
rect 2668 2076 2670 2079
rect 2626 2060 2628 2063
rect 2631 2060 2633 2062
rect 2652 2060 2654 2062
rect 2668 2060 2670 2072
rect 2684 2070 2686 2079
rect 2689 2077 2691 2079
rect 2684 2060 2686 2063
rect 2689 2060 2691 2062
rect 2705 2060 2707 2079
rect 2721 2076 2723 2079
rect 2726 2077 2728 2079
rect 2721 2060 2723 2072
rect 2726 2060 2728 2067
rect 2742 2060 2744 2079
rect 2758 2070 2760 2079
rect 2763 2077 2765 2079
rect 2784 2077 2786 2079
rect 2800 2076 2802 2079
rect 2758 2060 2760 2063
rect 2763 2060 2765 2062
rect 2784 2060 2786 2062
rect 2800 2060 2802 2072
rect 2816 2070 2818 2079
rect 2821 2077 2823 2079
rect 2837 2071 2839 2079
rect 2816 2060 2818 2063
rect 2821 2060 2823 2062
rect 2837 2060 2839 2067
rect 1512 2054 1514 2056
rect 1517 2053 1519 2056
rect 1533 2054 1535 2056
rect 1549 2054 1551 2056
rect 1554 2051 1556 2056
rect 1575 2051 1577 2056
rect 1591 2054 1593 2056
rect 1607 2054 1609 2056
rect 1612 2051 1614 2056
rect 1628 2054 1630 2056
rect 1644 2054 1646 2056
rect 1649 2053 1651 2056
rect 1665 2054 1667 2056
rect 1681 2054 1683 2056
rect 1686 2051 1688 2056
rect 1707 2051 1709 2056
rect 1723 2054 1725 2056
rect 1739 2054 1741 2056
rect 1744 2051 1746 2056
rect 1760 2054 1762 2056
rect 1776 2054 1778 2056
rect 1781 2053 1783 2056
rect 1797 2054 1799 2056
rect 1813 2054 1815 2056
rect 1818 2051 1820 2056
rect 1839 2051 1841 2056
rect 1855 2054 1857 2056
rect 1871 2054 1873 2056
rect 1876 2051 1878 2056
rect 1892 2054 1894 2056
rect 2457 2054 2459 2056
rect 2462 2053 2464 2056
rect 2478 2054 2480 2056
rect 2494 2054 2496 2056
rect 2499 2051 2501 2056
rect 2520 2051 2522 2056
rect 2536 2054 2538 2056
rect 2552 2054 2554 2056
rect 2557 2051 2559 2056
rect 2573 2054 2575 2056
rect 2589 2054 2591 2056
rect 2594 2053 2596 2056
rect 2610 2054 2612 2056
rect 2626 2054 2628 2056
rect 2631 2051 2633 2056
rect 2652 2051 2654 2056
rect 2668 2054 2670 2056
rect 2684 2054 2686 2056
rect 2689 2051 2691 2056
rect 2705 2054 2707 2056
rect 2721 2054 2723 2056
rect 2726 2053 2728 2056
rect 2742 2054 2744 2056
rect 2758 2054 2760 2056
rect 2763 2051 2765 2056
rect 2784 2051 2786 2056
rect 2800 2054 2802 2056
rect 2816 2054 2818 2056
rect 2821 2051 2823 2056
rect 2837 2054 2839 2056
rect 2295 2031 2297 2033
rect 2300 2031 2302 2034
rect 2316 2031 2318 2033
rect 2332 2031 2334 2033
rect 2337 2031 2339 2034
rect 2358 2031 2360 2034
rect 2374 2031 2376 2034
rect 2390 2031 2392 2033
rect 2395 2031 2397 2034
rect 2411 2031 2413 2033
rect 3240 2031 3242 2033
rect 3245 2031 3247 2034
rect 3261 2031 3263 2033
rect 3277 2031 3279 2033
rect 3282 2031 3284 2034
rect 3303 2031 3305 2034
rect 3319 2031 3321 2034
rect 3335 2031 3337 2033
rect 3340 2031 3342 2034
rect 3356 2031 3358 2033
rect 2295 2018 2297 2023
rect 2300 2021 2302 2023
rect 2295 2004 2297 2014
rect 2300 2004 2302 2011
rect 2316 2004 2318 2023
rect 2332 2014 2334 2023
rect 2337 2021 2339 2023
rect 2358 2021 2360 2023
rect 2374 2020 2376 2023
rect 2332 2004 2334 2007
rect 2337 2004 2339 2006
rect 2358 2004 2360 2006
rect 2374 2004 2376 2016
rect 2390 2014 2392 2023
rect 2395 2021 2397 2023
rect 2390 2004 2392 2007
rect 2395 2004 2397 2006
rect 2411 2004 2413 2023
rect 3240 2018 3242 2023
rect 3245 2021 3247 2023
rect 2433 2010 2436 2012
rect 2440 2010 2443 2012
rect 3240 2004 3242 2014
rect 3245 2004 3247 2011
rect 3261 2004 3263 2023
rect 3277 2014 3279 2023
rect 3282 2021 3284 2023
rect 3303 2021 3305 2023
rect 3319 2020 3321 2023
rect 3277 2004 3279 2007
rect 3282 2004 3284 2006
rect 3303 2004 3305 2006
rect 3319 2004 3321 2016
rect 3335 2014 3337 2023
rect 3340 2021 3342 2023
rect 3335 2004 3337 2007
rect 3340 2004 3342 2006
rect 3356 2004 3358 2023
rect 3378 2010 3381 2012
rect 3385 2010 3388 2012
rect 1512 2001 1514 2003
rect 1517 2001 1519 2004
rect 1533 2001 1535 2003
rect 1549 2001 1551 2003
rect 1554 2001 1556 2004
rect 1575 2001 1577 2004
rect 1591 2001 1593 2004
rect 1607 2001 1609 2003
rect 1612 2001 1614 2004
rect 1628 2001 1630 2003
rect 1644 2001 1646 2003
rect 1649 2001 1651 2004
rect 1665 2001 1667 2003
rect 1681 2001 1683 2003
rect 1686 2001 1688 2004
rect 1707 2001 1709 2004
rect 1723 2001 1725 2004
rect 1739 2001 1741 2003
rect 1744 2001 1746 2004
rect 1760 2001 1762 2003
rect 1776 2001 1778 2003
rect 1781 2001 1783 2004
rect 1797 2001 1799 2003
rect 1813 2001 1815 2003
rect 1818 2001 1820 2004
rect 1839 2001 1841 2004
rect 1855 2001 1857 2004
rect 1871 2001 1873 2003
rect 1876 2001 1878 2004
rect 1892 2001 1894 2003
rect 2457 2001 2459 2003
rect 2462 2001 2464 2004
rect 2478 2001 2480 2003
rect 2494 2001 2496 2003
rect 2499 2001 2501 2004
rect 2520 2001 2522 2004
rect 2536 2001 2538 2004
rect 2552 2001 2554 2003
rect 2557 2001 2559 2004
rect 2573 2001 2575 2003
rect 2589 2001 2591 2003
rect 2594 2001 2596 2004
rect 2610 2001 2612 2003
rect 2626 2001 2628 2003
rect 2631 2001 2633 2004
rect 2652 2001 2654 2004
rect 2668 2001 2670 2004
rect 2684 2001 2686 2003
rect 2689 2001 2691 2004
rect 2705 2001 2707 2003
rect 2721 2001 2723 2003
rect 2726 2001 2728 2004
rect 2742 2001 2744 2003
rect 2758 2001 2760 2003
rect 2763 2001 2765 2004
rect 2784 2001 2786 2004
rect 2800 2001 2802 2004
rect 2816 2001 2818 2003
rect 2821 2001 2823 2004
rect 2837 2001 2839 2003
rect 2295 1998 2297 2000
rect 2300 1997 2302 2000
rect 2316 1998 2318 2000
rect 2332 1998 2334 2000
rect 2337 1995 2339 2000
rect 2358 1995 2360 2000
rect 2374 1998 2376 2000
rect 2390 1998 2392 2000
rect 2395 1995 2397 2000
rect 2411 1998 2413 2000
rect 1512 1988 1514 1993
rect 1517 1991 1519 1993
rect 1512 1974 1514 1984
rect 1517 1974 1519 1981
rect 1533 1974 1535 1993
rect 1549 1984 1551 1993
rect 1554 1991 1556 1993
rect 1575 1991 1577 1993
rect 1591 1990 1593 1993
rect 1549 1974 1551 1977
rect 1554 1974 1556 1976
rect 1575 1974 1577 1976
rect 1591 1974 1593 1986
rect 1607 1984 1609 1993
rect 1612 1991 1614 1993
rect 1607 1974 1609 1977
rect 1612 1974 1614 1976
rect 1628 1974 1630 1993
rect 1644 1990 1646 1993
rect 1649 1991 1651 1993
rect 1644 1974 1646 1986
rect 1649 1974 1651 1981
rect 1665 1974 1667 1993
rect 1681 1984 1683 1993
rect 1686 1991 1688 1993
rect 1707 1991 1709 1993
rect 1723 1990 1725 1993
rect 1681 1974 1683 1977
rect 1686 1974 1688 1976
rect 1707 1974 1709 1976
rect 1723 1974 1725 1986
rect 1739 1984 1741 1993
rect 1744 1991 1746 1993
rect 1739 1974 1741 1977
rect 1744 1974 1746 1976
rect 1760 1974 1762 1993
rect 1776 1990 1778 1993
rect 1781 1991 1783 1993
rect 1776 1974 1778 1986
rect 1781 1974 1783 1981
rect 1797 1974 1799 1993
rect 1813 1984 1815 1993
rect 1818 1991 1820 1993
rect 1839 1991 1841 1993
rect 1855 1990 1857 1993
rect 1813 1974 1815 1977
rect 1818 1974 1820 1976
rect 1839 1974 1841 1976
rect 1855 1974 1857 1986
rect 1871 1984 1873 1993
rect 1876 1991 1878 1993
rect 1892 1985 1894 1993
rect 3240 1998 3242 2000
rect 3245 1997 3247 2000
rect 3261 1998 3263 2000
rect 3277 1998 3279 2000
rect 3282 1995 3284 2000
rect 3303 1995 3305 2000
rect 3319 1998 3321 2000
rect 3335 1998 3337 2000
rect 3340 1995 3342 2000
rect 3356 1998 3358 2000
rect 2457 1988 2459 1993
rect 2462 1991 2464 1993
rect 1871 1974 1873 1977
rect 1876 1974 1878 1976
rect 1892 1974 1894 1981
rect 2457 1974 2459 1984
rect 2462 1974 2464 1981
rect 2478 1974 2480 1993
rect 2494 1984 2496 1993
rect 2499 1991 2501 1993
rect 2520 1991 2522 1993
rect 2536 1990 2538 1993
rect 2494 1974 2496 1977
rect 2499 1974 2501 1976
rect 2520 1974 2522 1976
rect 2536 1974 2538 1986
rect 2552 1984 2554 1993
rect 2557 1991 2559 1993
rect 2552 1974 2554 1977
rect 2557 1974 2559 1976
rect 2573 1974 2575 1993
rect 2589 1990 2591 1993
rect 2594 1991 2596 1993
rect 2589 1974 2591 1986
rect 2594 1974 2596 1981
rect 2610 1974 2612 1993
rect 2626 1984 2628 1993
rect 2631 1991 2633 1993
rect 2652 1991 2654 1993
rect 2668 1990 2670 1993
rect 2626 1974 2628 1977
rect 2631 1974 2633 1976
rect 2652 1974 2654 1976
rect 2668 1974 2670 1986
rect 2684 1984 2686 1993
rect 2689 1991 2691 1993
rect 2684 1974 2686 1977
rect 2689 1974 2691 1976
rect 2705 1974 2707 1993
rect 2721 1990 2723 1993
rect 2726 1991 2728 1993
rect 2721 1974 2723 1986
rect 2726 1974 2728 1981
rect 2742 1974 2744 1993
rect 2758 1984 2760 1993
rect 2763 1991 2765 1993
rect 2784 1991 2786 1993
rect 2800 1990 2802 1993
rect 2758 1974 2760 1977
rect 2763 1974 2765 1976
rect 2784 1974 2786 1976
rect 2800 1974 2802 1986
rect 2816 1984 2818 1993
rect 2821 1991 2823 1993
rect 2837 1985 2839 1993
rect 2816 1974 2818 1977
rect 2821 1974 2823 1976
rect 2837 1974 2839 1981
rect 1512 1968 1514 1970
rect 1517 1967 1519 1970
rect 1533 1968 1535 1970
rect 1549 1968 1551 1970
rect 1554 1965 1556 1970
rect 1575 1965 1577 1970
rect 1591 1968 1593 1970
rect 1607 1968 1609 1970
rect 1612 1965 1614 1970
rect 1628 1968 1630 1970
rect 1644 1968 1646 1970
rect 1649 1967 1651 1970
rect 1665 1968 1667 1970
rect 1681 1968 1683 1970
rect 1686 1965 1688 1970
rect 1707 1965 1709 1970
rect 1723 1968 1725 1970
rect 1739 1968 1741 1970
rect 1744 1965 1746 1970
rect 1760 1968 1762 1970
rect 1776 1968 1778 1970
rect 1781 1967 1783 1970
rect 1797 1968 1799 1970
rect 1813 1968 1815 1970
rect 1818 1965 1820 1970
rect 1839 1965 1841 1970
rect 1855 1968 1857 1970
rect 1871 1968 1873 1970
rect 1876 1965 1878 1970
rect 1892 1968 1894 1970
rect 2457 1968 2459 1970
rect 2462 1967 2464 1970
rect 2478 1968 2480 1970
rect 2494 1968 2496 1970
rect 2499 1965 2501 1970
rect 2520 1965 2522 1970
rect 2536 1968 2538 1970
rect 2552 1968 2554 1970
rect 2557 1965 2559 1970
rect 2573 1968 2575 1970
rect 2589 1968 2591 1970
rect 2594 1967 2596 1970
rect 2610 1968 2612 1970
rect 2626 1968 2628 1970
rect 2631 1965 2633 1970
rect 2652 1965 2654 1970
rect 2668 1968 2670 1970
rect 2684 1968 2686 1970
rect 2689 1965 2691 1970
rect 2705 1968 2707 1970
rect 2721 1968 2723 1970
rect 2726 1967 2728 1970
rect 2742 1968 2744 1970
rect 2758 1968 2760 1970
rect 2763 1965 2765 1970
rect 2784 1965 2786 1970
rect 2800 1968 2802 1970
rect 2816 1968 2818 1970
rect 2821 1965 2823 1970
rect 2837 1968 2839 1970
rect 1744 1930 1746 1933
rect 1768 1930 1770 1933
rect 2689 1930 2691 1933
rect 2713 1930 2715 1933
rect 1744 1924 1746 1926
rect 1768 1924 1770 1926
rect 2689 1924 2691 1926
rect 2713 1924 2715 1926
rect 1764 1919 1766 1921
rect 2709 1919 2711 1921
rect 1764 1912 1766 1915
rect 2709 1912 2711 1915
rect 1753 1901 1755 1903
rect 1759 1901 1778 1903
rect 2698 1901 2700 1903
rect 2704 1901 2723 1903
rect 1744 1896 1746 1898
rect 1768 1896 1770 1898
rect 2689 1896 2691 1898
rect 2713 1896 2715 1898
rect 1744 1889 1746 1892
rect 1768 1889 1770 1892
rect 2689 1889 2691 1892
rect 2713 1889 2715 1892
rect 1512 1861 1514 1863
rect 1517 1861 1519 1864
rect 1533 1861 1535 1863
rect 1549 1861 1551 1863
rect 1554 1861 1556 1864
rect 1575 1861 1577 1864
rect 1591 1861 1593 1864
rect 1607 1861 1609 1863
rect 1612 1861 1614 1864
rect 1628 1861 1630 1863
rect 1644 1861 1646 1863
rect 1649 1861 1651 1864
rect 1665 1861 1667 1863
rect 1681 1861 1683 1863
rect 1686 1861 1688 1864
rect 1707 1861 1709 1864
rect 1723 1861 1725 1864
rect 1739 1861 1741 1863
rect 1744 1861 1746 1864
rect 1760 1861 1762 1863
rect 1776 1861 1778 1863
rect 1781 1861 1783 1864
rect 1797 1861 1799 1863
rect 1813 1861 1815 1863
rect 1818 1861 1820 1864
rect 1839 1861 1841 1864
rect 1855 1861 1857 1864
rect 1871 1861 1873 1863
rect 1876 1861 1878 1864
rect 1892 1861 1894 1863
rect 2457 1861 2459 1863
rect 2462 1861 2464 1864
rect 2478 1861 2480 1863
rect 2494 1861 2496 1863
rect 2499 1861 2501 1864
rect 2520 1861 2522 1864
rect 2536 1861 2538 1864
rect 2552 1861 2554 1863
rect 2557 1861 2559 1864
rect 2573 1861 2575 1863
rect 2589 1861 2591 1863
rect 2594 1861 2596 1864
rect 2610 1861 2612 1863
rect 2626 1861 2628 1863
rect 2631 1861 2633 1864
rect 2652 1861 2654 1864
rect 2668 1861 2670 1864
rect 2684 1861 2686 1863
rect 2689 1861 2691 1864
rect 2705 1861 2707 1863
rect 2721 1861 2723 1863
rect 2726 1861 2728 1864
rect 2742 1861 2744 1863
rect 2758 1861 2760 1863
rect 2763 1861 2765 1864
rect 2784 1861 2786 1864
rect 2800 1861 2802 1864
rect 2816 1861 2818 1863
rect 2821 1861 2823 1864
rect 2837 1861 2839 1863
rect 1512 1848 1514 1853
rect 1517 1851 1519 1853
rect 1512 1834 1514 1844
rect 1517 1834 1519 1841
rect 1533 1834 1535 1853
rect 1549 1844 1551 1853
rect 1554 1851 1556 1853
rect 1575 1851 1577 1853
rect 1591 1850 1593 1853
rect 1549 1834 1551 1837
rect 1554 1834 1556 1836
rect 1575 1834 1577 1836
rect 1591 1834 1593 1846
rect 1607 1844 1609 1853
rect 1612 1851 1614 1853
rect 1607 1834 1609 1837
rect 1612 1834 1614 1836
rect 1628 1834 1630 1853
rect 1644 1850 1646 1853
rect 1649 1851 1651 1853
rect 1644 1834 1646 1846
rect 1649 1834 1651 1841
rect 1665 1834 1667 1853
rect 1681 1844 1683 1853
rect 1686 1851 1688 1853
rect 1707 1851 1709 1853
rect 1723 1850 1725 1853
rect 1681 1834 1683 1837
rect 1686 1834 1688 1836
rect 1707 1834 1709 1836
rect 1723 1834 1725 1846
rect 1739 1844 1741 1853
rect 1744 1851 1746 1853
rect 1739 1834 1741 1837
rect 1744 1834 1746 1836
rect 1760 1834 1762 1853
rect 1776 1850 1778 1853
rect 1781 1851 1783 1853
rect 1776 1834 1778 1846
rect 1781 1834 1783 1841
rect 1797 1834 1799 1853
rect 1813 1844 1815 1853
rect 1818 1851 1820 1853
rect 1839 1851 1841 1853
rect 1855 1850 1857 1853
rect 1813 1834 1815 1837
rect 1818 1834 1820 1836
rect 1839 1834 1841 1836
rect 1855 1834 1857 1846
rect 1871 1844 1873 1853
rect 1876 1851 1878 1853
rect 1892 1845 1894 1853
rect 2457 1848 2459 1853
rect 2462 1851 2464 1853
rect 1871 1834 1873 1837
rect 1876 1834 1878 1836
rect 1892 1834 1894 1841
rect 2457 1834 2459 1844
rect 2462 1834 2464 1841
rect 2478 1834 2480 1853
rect 2494 1844 2496 1853
rect 2499 1851 2501 1853
rect 2520 1851 2522 1853
rect 2536 1850 2538 1853
rect 2494 1834 2496 1837
rect 2499 1834 2501 1836
rect 2520 1834 2522 1836
rect 2536 1834 2538 1846
rect 2552 1844 2554 1853
rect 2557 1851 2559 1853
rect 2552 1834 2554 1837
rect 2557 1834 2559 1836
rect 2573 1834 2575 1853
rect 2589 1850 2591 1853
rect 2594 1851 2596 1853
rect 2589 1834 2591 1846
rect 2594 1834 2596 1841
rect 2610 1834 2612 1853
rect 2626 1844 2628 1853
rect 2631 1851 2633 1853
rect 2652 1851 2654 1853
rect 2668 1850 2670 1853
rect 2626 1834 2628 1837
rect 2631 1834 2633 1836
rect 2652 1834 2654 1836
rect 2668 1834 2670 1846
rect 2684 1844 2686 1853
rect 2689 1851 2691 1853
rect 2684 1834 2686 1837
rect 2689 1834 2691 1836
rect 2705 1834 2707 1853
rect 2721 1850 2723 1853
rect 2726 1851 2728 1853
rect 2721 1834 2723 1846
rect 2726 1834 2728 1841
rect 2742 1834 2744 1853
rect 2758 1844 2760 1853
rect 2763 1851 2765 1853
rect 2784 1851 2786 1853
rect 2800 1850 2802 1853
rect 2758 1834 2760 1837
rect 2763 1834 2765 1836
rect 2784 1834 2786 1836
rect 2800 1834 2802 1846
rect 2816 1844 2818 1853
rect 2821 1851 2823 1853
rect 2837 1845 2839 1853
rect 2816 1834 2818 1837
rect 2821 1834 2823 1836
rect 2837 1834 2839 1841
rect 1512 1828 1514 1830
rect 1517 1827 1519 1830
rect 1533 1828 1535 1830
rect 1549 1828 1551 1830
rect 1554 1825 1556 1830
rect 1575 1825 1577 1830
rect 1591 1828 1593 1830
rect 1607 1828 1609 1830
rect 1612 1825 1614 1830
rect 1628 1828 1630 1830
rect 1644 1828 1646 1830
rect 1649 1827 1651 1830
rect 1665 1828 1667 1830
rect 1681 1828 1683 1830
rect 1686 1825 1688 1830
rect 1707 1825 1709 1830
rect 1723 1828 1725 1830
rect 1739 1828 1741 1830
rect 1744 1825 1746 1830
rect 1760 1828 1762 1830
rect 1776 1828 1778 1830
rect 1781 1827 1783 1830
rect 1797 1828 1799 1830
rect 1813 1828 1815 1830
rect 1818 1825 1820 1830
rect 1839 1825 1841 1830
rect 1855 1828 1857 1830
rect 1871 1828 1873 1830
rect 1876 1825 1878 1830
rect 1892 1828 1894 1830
rect 2457 1828 2459 1830
rect 2462 1827 2464 1830
rect 2478 1828 2480 1830
rect 2494 1828 2496 1830
rect 2499 1825 2501 1830
rect 2520 1825 2522 1830
rect 2536 1828 2538 1830
rect 2552 1828 2554 1830
rect 2557 1825 2559 1830
rect 2573 1828 2575 1830
rect 2589 1828 2591 1830
rect 2594 1827 2596 1830
rect 2610 1828 2612 1830
rect 2626 1828 2628 1830
rect 2631 1825 2633 1830
rect 2652 1825 2654 1830
rect 2668 1828 2670 1830
rect 2684 1828 2686 1830
rect 2689 1825 2691 1830
rect 2705 1828 2707 1830
rect 2721 1828 2723 1830
rect 2726 1827 2728 1830
rect 2742 1828 2744 1830
rect 2758 1828 2760 1830
rect 2763 1825 2765 1830
rect 2784 1825 2786 1830
rect 2800 1828 2802 1830
rect 2816 1828 2818 1830
rect 2821 1825 2823 1830
rect 2837 1828 2839 1830
<< polycontact >>
rect 2732 4273 2736 4277
rect 2697 4259 2701 4263
rect 2724 4255 2728 4259
rect 2751 4251 2755 4255
rect 2730 4237 2734 4241
rect 2885 4231 2889 4235
rect 2938 4231 2942 4235
rect 2732 4193 2736 4197
rect 2721 4177 2727 4181
rect 2730 4157 2734 4161
rect 2732 4143 2736 4147
rect 2675 4129 2679 4133
rect 2697 4129 2701 4133
rect 2724 4125 2728 4129
rect 2751 4121 2755 4125
rect 2730 4107 2734 4111
rect 2791 4101 2795 4105
rect 2844 4101 2848 4105
rect 2732 4063 2736 4067
rect 2721 4047 2727 4051
rect 2730 4027 2734 4031
rect 2001 3749 2005 3753
rect 2038 3749 2042 3753
rect 2058 3749 2062 3753
rect 2096 3749 2100 3753
rect 2133 3749 2137 3753
rect 2170 3749 2174 3753
rect 2190 3749 2194 3753
rect 2228 3749 2232 3753
rect 2265 3749 2269 3753
rect 2302 3749 2306 3753
rect 2322 3749 2326 3753
rect 2360 3749 2364 3753
rect 2397 3749 2401 3753
rect 2434 3749 2438 3753
rect 2454 3749 2458 3753
rect 2492 3749 2496 3753
rect 2946 3749 2950 3753
rect 2983 3749 2987 3753
rect 3003 3749 3007 3753
rect 3041 3749 3045 3753
rect 3078 3749 3082 3753
rect 3115 3749 3119 3753
rect 3135 3749 3139 3753
rect 3173 3749 3177 3753
rect 3210 3749 3214 3753
rect 3247 3749 3251 3753
rect 3267 3749 3271 3753
rect 3305 3749 3309 3753
rect 3342 3749 3346 3753
rect 3379 3749 3383 3753
rect 3399 3749 3403 3753
rect 3437 3749 3441 3753
rect 1995 3729 1999 3733
rect 2013 3731 2017 3735
rect 1649 3716 1653 3720
rect 1686 3716 1690 3720
rect 1706 3716 1710 3720
rect 1744 3716 1748 3720
rect 2073 3731 2077 3735
rect 2031 3722 2035 3729
rect 2089 3722 2093 3729
rect 2110 3726 2114 3730
rect 2127 3729 2131 3733
rect 2145 3731 2149 3735
rect 2205 3731 2209 3735
rect 2163 3722 2167 3729
rect 2221 3722 2225 3729
rect 2242 3726 2246 3730
rect 2259 3729 2263 3733
rect 2277 3731 2281 3735
rect 2337 3731 2341 3735
rect 2295 3722 2299 3729
rect 2353 3722 2357 3729
rect 2374 3726 2378 3730
rect 2391 3729 2395 3733
rect 2409 3731 2413 3735
rect 2469 3731 2473 3735
rect 2427 3722 2431 3729
rect 2485 3722 2489 3729
rect 2506 3726 2510 3730
rect 2940 3729 2944 3733
rect 2958 3731 2962 3735
rect 2594 3716 2598 3720
rect 2631 3716 2635 3720
rect 2651 3716 2655 3720
rect 2689 3716 2693 3720
rect 3018 3731 3022 3735
rect 2976 3722 2980 3729
rect 3034 3722 3038 3729
rect 3055 3726 3059 3730
rect 3072 3729 3076 3733
rect 3090 3731 3094 3735
rect 3150 3731 3154 3735
rect 3108 3722 3112 3729
rect 3166 3722 3170 3729
rect 3187 3726 3191 3730
rect 3204 3729 3208 3733
rect 3222 3731 3226 3735
rect 3282 3731 3286 3735
rect 3240 3722 3244 3729
rect 3298 3722 3302 3729
rect 3319 3726 3323 3730
rect 3336 3729 3340 3733
rect 3354 3731 3358 3735
rect 3414 3731 3418 3735
rect 3372 3722 3376 3729
rect 3430 3722 3434 3729
rect 3451 3726 3455 3730
rect 2001 3708 2005 3712
rect 2038 3706 2042 3710
rect 2058 3706 2062 3710
rect 2094 3706 2098 3710
rect 2133 3708 2137 3712
rect 2170 3706 2174 3710
rect 2190 3706 2194 3710
rect 2226 3706 2230 3710
rect 2265 3708 2269 3712
rect 2302 3706 2306 3710
rect 2322 3706 2326 3710
rect 2358 3706 2362 3710
rect 2397 3708 2401 3712
rect 2434 3706 2438 3710
rect 2454 3706 2458 3710
rect 2490 3706 2494 3710
rect 2946 3708 2950 3712
rect 2983 3706 2987 3710
rect 3003 3706 3007 3710
rect 3039 3706 3043 3710
rect 3078 3708 3082 3712
rect 3115 3706 3119 3710
rect 3135 3706 3139 3710
rect 3171 3706 3175 3710
rect 3210 3708 3214 3712
rect 3247 3706 3251 3710
rect 3267 3706 3271 3710
rect 3303 3706 3307 3710
rect 3342 3708 3346 3712
rect 3379 3706 3383 3710
rect 3399 3706 3403 3710
rect 3435 3706 3439 3710
rect 1643 3696 1647 3700
rect 1661 3698 1665 3702
rect 1721 3698 1725 3702
rect 1679 3689 1683 3696
rect 1737 3689 1741 3696
rect 1756 3693 1760 3697
rect 2588 3696 2592 3700
rect 2606 3698 2610 3702
rect 2666 3698 2670 3702
rect 2624 3689 2628 3696
rect 2682 3689 2686 3696
rect 2701 3693 2705 3697
rect 1649 3675 1653 3679
rect 1686 3673 1690 3677
rect 1706 3673 1710 3677
rect 1742 3673 1746 3677
rect 2017 3665 2021 3669
rect 2061 3665 2065 3669
rect 2088 3665 2092 3669
rect 2133 3665 2137 3669
rect 2206 3672 2210 3676
rect 1767 3652 1771 3656
rect 2171 3658 2175 3662
rect 1650 3643 1654 3647
rect 1997 3645 2001 3649
rect 2029 3646 2033 3650
rect 2048 3645 2052 3649
rect 2104 3646 2108 3650
rect 2120 3645 2124 3649
rect 2147 3645 2151 3649
rect 2287 3672 2291 3676
rect 2594 3675 2598 3679
rect 2198 3654 2202 3658
rect 2225 3650 2229 3654
rect 2252 3658 2256 3662
rect 2631 3673 2635 3677
rect 2651 3673 2655 3677
rect 2687 3673 2691 3677
rect 2279 3654 2283 3658
rect 2306 3650 2310 3654
rect 2962 3665 2966 3669
rect 3006 3665 3010 3669
rect 3033 3665 3037 3669
rect 3078 3665 3082 3669
rect 3151 3672 3155 3676
rect 2712 3652 2716 3656
rect 3116 3658 3120 3662
rect 2204 3636 2208 3640
rect 2595 3643 2599 3647
rect 2942 3645 2946 3649
rect 2285 3636 2289 3640
rect 2974 3646 2978 3650
rect 2993 3645 2997 3649
rect 3049 3646 3053 3650
rect 3065 3645 3069 3649
rect 3092 3645 3096 3649
rect 3232 3672 3236 3676
rect 3143 3654 3147 3658
rect 3170 3650 3174 3654
rect 3197 3658 3201 3662
rect 3224 3654 3228 3658
rect 3251 3650 3255 3654
rect 3149 3636 3153 3640
rect 3230 3636 3234 3640
rect 2014 3628 2018 3632
rect 2058 3627 2062 3631
rect 2083 3628 2088 3632
rect 2130 3627 2134 3631
rect 2959 3628 2963 3632
rect 3003 3627 3007 3631
rect 3028 3628 3033 3632
rect 3075 3627 3079 3631
rect 1649 3614 1653 3618
rect 1687 3614 1691 3618
rect 1707 3614 1711 3618
rect 1744 3614 1748 3618
rect 2594 3614 2598 3618
rect 2632 3614 2636 3618
rect 2652 3614 2656 3618
rect 2689 3614 2693 3618
rect 1637 3591 1641 3595
rect 1672 3596 1676 3600
rect 1656 3587 1660 3594
rect 1714 3587 1718 3594
rect 1732 3596 1736 3600
rect 2014 3598 2018 3602
rect 2058 3599 2062 3603
rect 1750 3594 1754 3598
rect 2083 3598 2088 3602
rect 2130 3599 2134 3603
rect 2206 3596 2210 3600
rect 2287 3596 2291 3600
rect 1997 3581 2001 3585
rect 1651 3571 1655 3575
rect 1687 3571 1691 3575
rect 1707 3571 1711 3575
rect 1744 3573 1748 3577
rect 2029 3580 2033 3584
rect 2048 3581 2052 3585
rect 2104 3580 2108 3584
rect 2120 3581 2124 3585
rect 2147 3581 2151 3585
rect 2195 3580 2201 3584
rect 2276 3580 2282 3584
rect 2582 3591 2586 3595
rect 2617 3596 2621 3600
rect 2601 3587 2605 3594
rect 2659 3587 2663 3594
rect 2677 3596 2681 3600
rect 2959 3598 2963 3602
rect 3003 3599 3007 3603
rect 2695 3594 2699 3598
rect 3028 3598 3033 3602
rect 3075 3599 3079 3603
rect 3151 3596 3155 3600
rect 3232 3596 3236 3600
rect 2942 3581 2946 3585
rect 2596 3571 2600 3575
rect 2632 3571 2636 3575
rect 2652 3571 2656 3575
rect 2689 3573 2693 3577
rect 2974 3580 2978 3584
rect 2993 3581 2997 3585
rect 3049 3580 3053 3584
rect 3065 3581 3069 3585
rect 3092 3581 3096 3585
rect 3140 3580 3146 3584
rect 3221 3580 3227 3584
rect 2017 3561 2021 3565
rect 2061 3561 2065 3565
rect 2088 3561 2092 3565
rect 2133 3561 2137 3565
rect 2204 3560 2208 3564
rect 2285 3560 2289 3564
rect 2962 3561 2966 3565
rect 3006 3561 3010 3565
rect 3033 3561 3037 3565
rect 3078 3561 3082 3565
rect 3149 3560 3153 3564
rect 3230 3560 3234 3564
rect 2206 3540 2210 3544
rect 2017 3533 2021 3537
rect 2061 3533 2065 3537
rect 2088 3533 2092 3537
rect 2133 3533 2137 3537
rect 2311 3540 2315 3544
rect 2198 3522 2202 3526
rect 1997 3513 2001 3517
rect 2029 3514 2033 3518
rect 2048 3513 2052 3517
rect 2104 3514 2108 3518
rect 2120 3513 2124 3517
rect 2147 3513 2151 3517
rect 2225 3518 2229 3522
rect 2276 3526 2280 3530
rect 3151 3540 3155 3544
rect 2303 3522 2307 3526
rect 2330 3518 2334 3522
rect 2962 3533 2966 3537
rect 3006 3533 3010 3537
rect 3033 3533 3037 3537
rect 3078 3533 3082 3537
rect 3256 3540 3260 3544
rect 3143 3522 3147 3526
rect 2942 3513 2946 3517
rect 2204 3504 2208 3508
rect 2309 3504 2313 3508
rect 2974 3514 2978 3518
rect 2993 3513 2997 3517
rect 3049 3514 3053 3518
rect 3065 3513 3069 3517
rect 3092 3513 3096 3517
rect 3170 3518 3174 3522
rect 3221 3526 3225 3530
rect 3248 3522 3252 3526
rect 3275 3518 3279 3522
rect 3149 3504 3153 3508
rect 3254 3504 3258 3508
rect 2014 3496 2018 3500
rect 2058 3495 2062 3499
rect 2083 3496 2088 3500
rect 2130 3495 2134 3499
rect 2959 3496 2963 3500
rect 3003 3495 3007 3499
rect 3028 3496 3033 3500
rect 3075 3495 3079 3499
rect 2014 3466 2018 3470
rect 2058 3467 2062 3471
rect 2083 3466 2088 3470
rect 2130 3467 2134 3471
rect 2206 3465 2210 3469
rect 2311 3465 2315 3469
rect 2959 3466 2963 3470
rect 3003 3467 3007 3471
rect 3028 3466 3033 3470
rect 3075 3467 3079 3471
rect 3151 3465 3155 3469
rect 3256 3465 3260 3469
rect 1997 3449 2001 3453
rect 2029 3448 2033 3452
rect 2048 3449 2052 3453
rect 2104 3448 2108 3452
rect 2120 3449 2124 3453
rect 2147 3449 2151 3453
rect 2195 3449 2201 3453
rect 2300 3449 2306 3453
rect 2942 3449 2946 3453
rect 2974 3448 2978 3452
rect 2993 3449 2997 3453
rect 3049 3448 3053 3452
rect 3065 3449 3069 3453
rect 3092 3449 3096 3453
rect 3140 3449 3146 3453
rect 3245 3449 3251 3453
rect 2017 3429 2021 3433
rect 2061 3429 2065 3433
rect 2088 3429 2092 3433
rect 2133 3429 2137 3433
rect 2204 3429 2208 3433
rect 2309 3429 2313 3433
rect 2962 3429 2966 3433
rect 3006 3429 3010 3433
rect 3033 3429 3037 3433
rect 3078 3429 3082 3433
rect 3149 3429 3153 3433
rect 3254 3429 3258 3433
rect 2206 3408 2210 3412
rect 2017 3401 2021 3405
rect 2061 3401 2065 3405
rect 2088 3401 2092 3405
rect 2133 3401 2137 3405
rect 2287 3408 2291 3412
rect 2198 3390 2202 3394
rect 1997 3381 2001 3385
rect 2029 3382 2033 3386
rect 2048 3381 2052 3385
rect 2104 3382 2108 3386
rect 2120 3381 2124 3385
rect 2147 3381 2151 3385
rect 2225 3386 2229 3390
rect 2252 3394 2256 3398
rect 2377 3408 2381 3412
rect 2279 3390 2283 3394
rect 2306 3386 2310 3390
rect 2342 3394 2346 3398
rect 3151 3408 3155 3412
rect 2369 3390 2373 3394
rect 2396 3386 2400 3390
rect 2962 3401 2966 3405
rect 3006 3401 3010 3405
rect 3033 3401 3037 3405
rect 3078 3401 3082 3405
rect 3232 3408 3236 3412
rect 3143 3390 3147 3394
rect 2942 3381 2946 3385
rect 2204 3372 2208 3376
rect 2285 3372 2289 3376
rect 2375 3372 2379 3376
rect 2974 3382 2978 3386
rect 2993 3381 2997 3385
rect 3049 3382 3053 3386
rect 3065 3381 3069 3385
rect 3092 3381 3096 3385
rect 3170 3386 3174 3390
rect 3197 3394 3201 3398
rect 3322 3408 3326 3412
rect 3224 3390 3228 3394
rect 3251 3386 3255 3390
rect 3287 3394 3291 3398
rect 3314 3390 3318 3394
rect 3341 3386 3345 3390
rect 3149 3372 3153 3376
rect 3230 3372 3234 3376
rect 3320 3372 3324 3376
rect 2014 3364 2018 3368
rect 2058 3363 2062 3367
rect 2083 3364 2088 3368
rect 2130 3363 2134 3367
rect 2959 3364 2963 3368
rect 3003 3363 3007 3367
rect 3028 3364 3033 3368
rect 3075 3363 3079 3367
rect 2014 3334 2018 3338
rect 2058 3335 2062 3339
rect 2083 3334 2088 3338
rect 2130 3335 2134 3339
rect 2959 3334 2963 3338
rect 3003 3335 3007 3339
rect 2206 3330 2210 3334
rect 2287 3330 2291 3334
rect 2377 3330 2381 3334
rect 3028 3334 3033 3338
rect 3075 3335 3079 3339
rect 3151 3330 3155 3334
rect 3232 3330 3236 3334
rect 3322 3330 3326 3334
rect 1997 3317 2001 3321
rect 2029 3316 2033 3320
rect 2048 3317 2052 3321
rect 2104 3316 2108 3320
rect 2120 3317 2124 3321
rect 2147 3317 2151 3321
rect 2195 3314 2201 3318
rect 2276 3314 2282 3318
rect 2366 3314 2372 3318
rect 2942 3317 2946 3321
rect 2974 3316 2978 3320
rect 2993 3317 2997 3321
rect 3049 3316 3053 3320
rect 3065 3317 3069 3321
rect 3092 3317 3096 3321
rect 3140 3314 3146 3318
rect 3221 3314 3227 3318
rect 3311 3314 3317 3318
rect 2017 3297 2021 3301
rect 2061 3297 2065 3301
rect 2088 3297 2092 3301
rect 2133 3297 2137 3301
rect 2204 3294 2208 3298
rect 2285 3294 2289 3298
rect 2375 3294 2379 3298
rect 2962 3297 2966 3301
rect 3006 3297 3010 3301
rect 3033 3297 3037 3301
rect 3078 3297 3082 3301
rect 3149 3294 3153 3298
rect 3230 3294 3234 3298
rect 3320 3294 3324 3298
rect 2206 3276 2210 3280
rect 2017 3269 2021 3273
rect 2061 3269 2065 3273
rect 2088 3269 2092 3273
rect 2133 3269 2137 3273
rect 3151 3276 3155 3280
rect 2198 3258 2202 3262
rect 1997 3249 2001 3253
rect 2029 3250 2033 3254
rect 2048 3249 2052 3253
rect 2104 3250 2108 3254
rect 2120 3249 2124 3253
rect 2147 3249 2151 3253
rect 2225 3254 2229 3258
rect 2962 3269 2966 3273
rect 3006 3269 3010 3273
rect 3033 3269 3037 3273
rect 3078 3269 3082 3273
rect 3143 3258 3147 3262
rect 2942 3249 2946 3253
rect 2204 3240 2208 3244
rect 2974 3250 2978 3254
rect 2993 3249 2997 3253
rect 3049 3250 3053 3254
rect 3065 3249 3069 3253
rect 3092 3249 3096 3253
rect 3170 3254 3174 3258
rect 3149 3240 3153 3244
rect 2014 3232 2018 3236
rect 2058 3231 2062 3235
rect 2083 3232 2088 3236
rect 2130 3231 2134 3235
rect 2959 3232 2963 3236
rect 3003 3231 3007 3235
rect 3028 3232 3033 3236
rect 3075 3231 3079 3235
rect 1517 3214 1521 3218
rect 1554 3214 1558 3218
rect 1574 3214 1578 3218
rect 1612 3214 1616 3218
rect 1649 3214 1653 3218
rect 1686 3214 1690 3218
rect 1706 3214 1710 3218
rect 1744 3214 1748 3218
rect 1781 3214 1785 3218
rect 1818 3214 1822 3218
rect 1838 3214 1842 3218
rect 1876 3214 1880 3218
rect 2462 3214 2466 3218
rect 2499 3214 2503 3218
rect 2519 3214 2523 3218
rect 2557 3214 2561 3218
rect 2594 3214 2598 3218
rect 2631 3214 2635 3218
rect 2651 3214 2655 3218
rect 2689 3214 2693 3218
rect 2726 3214 2730 3218
rect 2763 3214 2767 3218
rect 2783 3214 2787 3218
rect 2821 3214 2825 3218
rect 1511 3194 1515 3198
rect 1529 3196 1533 3200
rect 1589 3196 1593 3200
rect 1547 3187 1551 3194
rect 1605 3187 1609 3194
rect 1624 3191 1628 3195
rect 1642 3196 1646 3200
rect 1661 3196 1665 3200
rect 1721 3196 1725 3200
rect 1679 3187 1683 3194
rect 1737 3187 1741 3194
rect 1756 3191 1760 3195
rect 1774 3196 1778 3200
rect 1793 3196 1797 3200
rect 1853 3196 1857 3200
rect 1811 3187 1815 3194
rect 2014 3202 2018 3206
rect 2058 3203 2062 3207
rect 2083 3202 2088 3206
rect 2130 3203 2134 3207
rect 2275 3202 2279 3206
rect 2319 3203 2323 3207
rect 2344 3202 2349 3206
rect 2391 3203 2395 3207
rect 1869 3187 1873 3194
rect 1890 3191 1894 3195
rect 2206 3194 2210 3198
rect 2456 3194 2460 3198
rect 2474 3196 2478 3200
rect 1997 3185 2001 3189
rect 2029 3184 2033 3188
rect 2048 3185 2052 3189
rect 2104 3184 2108 3188
rect 2120 3185 2124 3189
rect 2147 3185 2151 3189
rect 1517 3173 1521 3177
rect 1554 3171 1558 3175
rect 1574 3171 1578 3175
rect 1610 3171 1614 3175
rect 1649 3173 1653 3177
rect 1686 3171 1690 3175
rect 1706 3171 1710 3175
rect 1742 3171 1746 3175
rect 1781 3173 1785 3177
rect 1818 3171 1822 3175
rect 1838 3171 1842 3175
rect 1874 3171 1878 3175
rect 2195 3178 2201 3182
rect 2233 3185 2237 3189
rect 2290 3184 2294 3188
rect 2309 3185 2313 3189
rect 2365 3184 2369 3188
rect 2381 3185 2385 3189
rect 2408 3185 2412 3189
rect 2534 3196 2538 3200
rect 2492 3187 2496 3194
rect 2550 3187 2554 3194
rect 2569 3191 2573 3195
rect 2587 3196 2591 3200
rect 2606 3196 2610 3200
rect 2666 3196 2670 3200
rect 2624 3187 2628 3194
rect 2682 3187 2686 3194
rect 2701 3191 2705 3195
rect 2719 3196 2723 3200
rect 2738 3196 2742 3200
rect 2798 3196 2802 3200
rect 2756 3187 2760 3194
rect 2959 3202 2963 3206
rect 3003 3203 3007 3207
rect 3028 3202 3033 3206
rect 3075 3203 3079 3207
rect 3220 3202 3224 3206
rect 3264 3203 3268 3207
rect 3289 3202 3294 3206
rect 3336 3203 3340 3207
rect 2814 3187 2818 3194
rect 2835 3191 2839 3195
rect 3151 3194 3155 3198
rect 2942 3185 2946 3189
rect 2974 3184 2978 3188
rect 2993 3185 2997 3189
rect 3049 3184 3053 3188
rect 3065 3185 3069 3189
rect 3092 3185 3096 3189
rect 2017 3165 2021 3169
rect 2061 3165 2065 3169
rect 2088 3165 2092 3169
rect 2133 3165 2137 3169
rect 2462 3173 2466 3177
rect 2204 3158 2208 3162
rect 1626 3143 1630 3147
rect 1650 3143 1654 3147
rect 2499 3171 2503 3175
rect 2519 3171 2523 3175
rect 2555 3171 2559 3175
rect 2594 3173 2598 3177
rect 2631 3171 2635 3175
rect 2651 3171 2655 3175
rect 2687 3171 2691 3175
rect 2726 3173 2730 3177
rect 2763 3171 2767 3175
rect 2783 3171 2787 3175
rect 2819 3171 2823 3175
rect 3140 3178 3146 3182
rect 3178 3185 3182 3189
rect 3235 3184 3239 3188
rect 3254 3185 3258 3189
rect 3310 3184 3314 3188
rect 3326 3185 3330 3189
rect 3353 3185 3357 3189
rect 2278 3165 2282 3169
rect 2322 3165 2326 3169
rect 2349 3165 2353 3169
rect 2394 3165 2398 3169
rect 2962 3165 2966 3169
rect 3006 3165 3010 3169
rect 3033 3165 3037 3169
rect 3078 3165 3082 3169
rect 3149 3158 3153 3162
rect 2571 3143 2575 3147
rect 2595 3143 2599 3147
rect 2417 3137 2421 3141
rect 2255 3130 2259 3134
rect 3223 3165 3227 3169
rect 3267 3165 3271 3169
rect 3294 3165 3298 3169
rect 3339 3165 3343 3169
rect 3362 3137 3366 3141
rect 3198 3130 3202 3134
rect 1646 3116 1650 3120
rect 2591 3116 2595 3120
rect 1661 3108 1665 3112
rect 2606 3108 2610 3112
rect 2300 3102 2304 3106
rect 2337 3102 2341 3106
rect 2357 3102 2361 3106
rect 2395 3102 2399 3106
rect 3245 3102 3249 3106
rect 3282 3102 3286 3106
rect 3302 3102 3306 3106
rect 3340 3102 3344 3106
rect 1626 3093 1630 3097
rect 1650 3093 1654 3097
rect 2571 3093 2575 3097
rect 2595 3093 2599 3097
rect 2294 3082 2298 3086
rect 2312 3084 2316 3088
rect 1517 3072 1521 3076
rect 1554 3072 1558 3076
rect 1574 3072 1578 3076
rect 1612 3072 1616 3076
rect 1649 3072 1653 3076
rect 1686 3072 1690 3076
rect 1706 3072 1710 3076
rect 1744 3072 1748 3076
rect 1781 3072 1785 3076
rect 1818 3072 1822 3076
rect 1838 3072 1842 3076
rect 1876 3072 1880 3076
rect 2372 3084 2376 3088
rect 2330 3075 2334 3082
rect 2388 3075 2392 3082
rect 2407 3079 2411 3083
rect 3239 3082 3243 3086
rect 3257 3084 3261 3088
rect 2462 3072 2466 3076
rect 2499 3072 2503 3076
rect 2519 3072 2523 3076
rect 2557 3072 2561 3076
rect 2594 3072 2598 3076
rect 2631 3072 2635 3076
rect 2651 3072 2655 3076
rect 2689 3072 2693 3076
rect 2726 3072 2730 3076
rect 2763 3072 2767 3076
rect 2783 3072 2787 3076
rect 2821 3072 2825 3076
rect 3317 3084 3321 3088
rect 3275 3075 3279 3082
rect 3333 3075 3337 3082
rect 3352 3079 3356 3083
rect 2300 3061 2304 3065
rect 1511 3052 1515 3056
rect 1529 3054 1533 3058
rect 1589 3054 1593 3058
rect 1547 3045 1551 3052
rect 1605 3045 1609 3052
rect 1624 3049 1628 3053
rect 1642 3054 1646 3058
rect 1661 3054 1665 3058
rect 1721 3054 1725 3058
rect 1679 3045 1683 3052
rect 1737 3045 1741 3052
rect 1756 3049 1760 3053
rect 1774 3054 1778 3058
rect 1793 3054 1797 3058
rect 1853 3054 1857 3058
rect 1811 3045 1815 3052
rect 2337 3059 2341 3063
rect 2357 3059 2361 3063
rect 2393 3059 2397 3063
rect 3245 3061 3249 3065
rect 1869 3045 1873 3052
rect 1890 3049 1894 3053
rect 2456 3052 2460 3056
rect 2474 3054 2478 3058
rect 2534 3054 2538 3058
rect 2492 3045 2496 3052
rect 2550 3045 2554 3052
rect 2569 3049 2573 3053
rect 2587 3054 2591 3058
rect 2606 3054 2610 3058
rect 2666 3054 2670 3058
rect 2624 3045 2628 3052
rect 2682 3045 2686 3052
rect 2701 3049 2705 3053
rect 2719 3054 2723 3058
rect 2738 3054 2742 3058
rect 2798 3054 2802 3058
rect 2756 3045 2760 3052
rect 3282 3059 3286 3063
rect 3302 3059 3306 3063
rect 3338 3059 3342 3063
rect 2814 3045 2818 3052
rect 2835 3049 2839 3053
rect 1517 3031 1521 3035
rect 1554 3029 1558 3033
rect 1574 3029 1578 3033
rect 1610 3029 1614 3033
rect 1649 3031 1653 3035
rect 1686 3029 1690 3033
rect 1706 3029 1710 3033
rect 1742 3029 1746 3033
rect 1781 3031 1785 3035
rect 1818 3029 1822 3033
rect 1838 3029 1842 3033
rect 1874 3029 1878 3033
rect 2462 3031 2466 3035
rect 2499 3029 2503 3033
rect 2519 3029 2523 3033
rect 2555 3029 2559 3033
rect 2594 3031 2598 3035
rect 2631 3029 2635 3033
rect 2651 3029 2655 3033
rect 2687 3029 2691 3033
rect 2726 3031 2730 3035
rect 2763 3029 2767 3033
rect 2783 3029 2787 3033
rect 2819 3029 2823 3033
rect 2300 3016 2304 3020
rect 2337 3016 2341 3020
rect 2357 3016 2361 3020
rect 2395 3016 2399 3020
rect 3245 3016 3249 3020
rect 3282 3016 3286 3020
rect 3302 3016 3306 3020
rect 3340 3016 3344 3020
rect 2294 2996 2298 3000
rect 2312 2998 2316 3002
rect 1517 2986 1521 2990
rect 1554 2986 1558 2990
rect 1574 2986 1578 2990
rect 1612 2986 1616 2990
rect 1649 2986 1653 2990
rect 1686 2986 1690 2990
rect 1706 2986 1710 2990
rect 1744 2986 1748 2990
rect 1781 2986 1785 2990
rect 1818 2986 1822 2990
rect 1838 2986 1842 2990
rect 1876 2986 1880 2990
rect 2372 2998 2376 3002
rect 2330 2989 2334 2996
rect 2388 2989 2392 2996
rect 2407 2993 2411 2997
rect 2429 2991 2433 2995
rect 3239 2996 3243 3000
rect 3257 2998 3261 3002
rect 2462 2986 2466 2990
rect 2499 2986 2503 2990
rect 2519 2986 2523 2990
rect 2557 2986 2561 2990
rect 2594 2986 2598 2990
rect 2631 2986 2635 2990
rect 2651 2986 2655 2990
rect 2689 2986 2693 2990
rect 2726 2986 2730 2990
rect 2763 2986 2767 2990
rect 2783 2986 2787 2990
rect 2821 2986 2825 2990
rect 3317 2998 3321 3002
rect 3275 2989 3279 2996
rect 3333 2989 3337 2996
rect 3352 2993 3356 2997
rect 3374 2991 3378 2995
rect 2300 2975 2304 2979
rect 1511 2966 1515 2970
rect 1529 2968 1533 2972
rect 1589 2968 1593 2972
rect 1547 2959 1551 2966
rect 1605 2959 1609 2966
rect 1624 2963 1628 2967
rect 1642 2968 1646 2972
rect 1661 2968 1665 2972
rect 1721 2968 1725 2972
rect 1679 2959 1683 2966
rect 1737 2959 1741 2966
rect 1756 2963 1760 2967
rect 1774 2968 1778 2972
rect 1793 2968 1797 2972
rect 1853 2968 1857 2972
rect 1811 2959 1815 2966
rect 2337 2973 2341 2977
rect 2357 2973 2361 2977
rect 2393 2973 2397 2977
rect 3245 2975 3249 2979
rect 1869 2959 1873 2966
rect 1890 2963 1894 2967
rect 2456 2966 2460 2970
rect 2474 2968 2478 2972
rect 2534 2968 2538 2972
rect 2492 2959 2496 2966
rect 2550 2959 2554 2966
rect 2569 2963 2573 2967
rect 2587 2968 2591 2972
rect 2606 2968 2610 2972
rect 2666 2968 2670 2972
rect 2624 2959 2628 2966
rect 2682 2959 2686 2966
rect 2701 2963 2705 2967
rect 2719 2968 2723 2972
rect 2738 2968 2742 2972
rect 2798 2968 2802 2972
rect 2756 2959 2760 2966
rect 3282 2973 3286 2977
rect 3302 2973 3306 2977
rect 3338 2973 3342 2977
rect 2814 2959 2818 2966
rect 2835 2963 2839 2967
rect 1517 2945 1521 2949
rect 1554 2943 1558 2947
rect 1574 2943 1578 2947
rect 1610 2943 1614 2947
rect 1649 2945 1653 2949
rect 1686 2943 1690 2947
rect 1706 2943 1710 2947
rect 1742 2943 1746 2947
rect 1781 2945 1785 2949
rect 1818 2943 1822 2947
rect 1838 2943 1842 2947
rect 1874 2943 1878 2947
rect 2462 2945 2466 2949
rect 2499 2943 2503 2947
rect 2519 2943 2523 2947
rect 2555 2943 2559 2947
rect 2594 2945 2598 2949
rect 2631 2943 2635 2947
rect 2651 2943 2655 2947
rect 2687 2943 2691 2947
rect 2726 2945 2730 2949
rect 2763 2943 2767 2947
rect 2783 2943 2787 2947
rect 2819 2943 2823 2947
rect 1743 2915 1747 2919
rect 1767 2915 1771 2919
rect 2688 2915 2692 2919
rect 2712 2915 2716 2919
rect 1763 2890 1767 2894
rect 2708 2890 2712 2894
rect 1778 2882 1782 2886
rect 2723 2882 2727 2886
rect 1743 2867 1747 2871
rect 1767 2867 1771 2871
rect 2688 2867 2692 2871
rect 2712 2867 2716 2871
rect 1517 2846 1521 2850
rect 1554 2846 1558 2850
rect 1574 2846 1578 2850
rect 1612 2846 1616 2850
rect 1649 2846 1653 2850
rect 1686 2846 1690 2850
rect 1706 2846 1710 2850
rect 1744 2846 1748 2850
rect 1781 2846 1785 2850
rect 1818 2846 1822 2850
rect 1838 2846 1842 2850
rect 1876 2846 1880 2850
rect 2462 2846 2466 2850
rect 2499 2846 2503 2850
rect 2519 2846 2523 2850
rect 2557 2846 2561 2850
rect 2594 2846 2598 2850
rect 2631 2846 2635 2850
rect 2651 2846 2655 2850
rect 2689 2846 2693 2850
rect 2726 2846 2730 2850
rect 2763 2846 2767 2850
rect 2783 2846 2787 2850
rect 2821 2846 2825 2850
rect 1511 2826 1515 2830
rect 1529 2828 1533 2832
rect 1589 2828 1593 2832
rect 1547 2819 1551 2826
rect 1605 2819 1609 2826
rect 1624 2823 1628 2827
rect 1642 2828 1646 2832
rect 1661 2828 1665 2832
rect 1721 2828 1725 2832
rect 1679 2819 1683 2826
rect 1737 2819 1741 2826
rect 1756 2823 1760 2827
rect 1774 2828 1778 2832
rect 1793 2828 1797 2832
rect 1853 2828 1857 2832
rect 1811 2819 1815 2826
rect 1869 2819 1873 2826
rect 1890 2823 1894 2827
rect 2456 2826 2460 2830
rect 2474 2828 2478 2832
rect 2534 2828 2538 2832
rect 2492 2819 2496 2826
rect 2550 2819 2554 2826
rect 2569 2823 2573 2827
rect 2587 2828 2591 2832
rect 2606 2828 2610 2832
rect 2666 2828 2670 2832
rect 2624 2819 2628 2826
rect 2682 2819 2686 2826
rect 2701 2823 2705 2827
rect 2719 2828 2723 2832
rect 2738 2828 2742 2832
rect 2798 2828 2802 2832
rect 2756 2819 2760 2826
rect 2814 2819 2818 2826
rect 2835 2823 2839 2827
rect 1517 2805 1521 2809
rect 1554 2803 1558 2807
rect 1574 2803 1578 2807
rect 1610 2803 1614 2807
rect 1649 2805 1653 2809
rect 1686 2803 1690 2807
rect 1706 2803 1710 2807
rect 1742 2803 1746 2807
rect 1781 2805 1785 2809
rect 1818 2803 1822 2807
rect 1838 2803 1842 2807
rect 1874 2803 1878 2807
rect 2462 2805 2466 2809
rect 2499 2803 2503 2807
rect 2519 2803 2523 2807
rect 2555 2803 2559 2807
rect 2594 2805 2598 2809
rect 2631 2803 2635 2807
rect 2651 2803 2655 2807
rect 2687 2803 2691 2807
rect 2726 2805 2730 2809
rect 2763 2803 2767 2807
rect 2783 2803 2787 2807
rect 2819 2803 2823 2807
rect 2001 2767 2005 2771
rect 2038 2767 2042 2771
rect 2058 2767 2062 2771
rect 2096 2767 2100 2771
rect 2133 2767 2137 2771
rect 2170 2767 2174 2771
rect 2190 2767 2194 2771
rect 2228 2767 2232 2771
rect 2265 2767 2269 2771
rect 2302 2767 2306 2771
rect 2322 2767 2326 2771
rect 2360 2767 2364 2771
rect 2397 2767 2401 2771
rect 2434 2767 2438 2771
rect 2454 2767 2458 2771
rect 2492 2767 2496 2771
rect 2946 2767 2950 2771
rect 2983 2767 2987 2771
rect 3003 2767 3007 2771
rect 3041 2767 3045 2771
rect 3078 2767 3082 2771
rect 3115 2767 3119 2771
rect 3135 2767 3139 2771
rect 3173 2767 3177 2771
rect 3210 2767 3214 2771
rect 3247 2767 3251 2771
rect 3267 2767 3271 2771
rect 3305 2767 3309 2771
rect 3342 2767 3346 2771
rect 3379 2767 3383 2771
rect 3399 2767 3403 2771
rect 3437 2767 3441 2771
rect 1995 2747 1999 2751
rect 2013 2749 2017 2753
rect 1649 2734 1653 2738
rect 1686 2734 1690 2738
rect 1706 2734 1710 2738
rect 1744 2734 1748 2738
rect 2073 2749 2077 2753
rect 2031 2740 2035 2747
rect 2089 2740 2093 2747
rect 2110 2744 2114 2748
rect 2127 2747 2131 2751
rect 2145 2749 2149 2753
rect 2205 2749 2209 2753
rect 2163 2740 2167 2747
rect 2221 2740 2225 2747
rect 2242 2744 2246 2748
rect 2259 2747 2263 2751
rect 2277 2749 2281 2753
rect 2337 2749 2341 2753
rect 2295 2740 2299 2747
rect 2353 2740 2357 2747
rect 2374 2744 2378 2748
rect 2391 2747 2395 2751
rect 2409 2749 2413 2753
rect 2469 2749 2473 2753
rect 2427 2740 2431 2747
rect 2485 2740 2489 2747
rect 2506 2744 2510 2748
rect 2940 2747 2944 2751
rect 2958 2749 2962 2753
rect 2594 2734 2598 2738
rect 2631 2734 2635 2738
rect 2651 2734 2655 2738
rect 2689 2734 2693 2738
rect 3018 2749 3022 2753
rect 2976 2740 2980 2747
rect 3034 2740 3038 2747
rect 3055 2744 3059 2748
rect 3072 2747 3076 2751
rect 3090 2749 3094 2753
rect 3150 2749 3154 2753
rect 3108 2740 3112 2747
rect 3166 2740 3170 2747
rect 3187 2744 3191 2748
rect 3204 2747 3208 2751
rect 3222 2749 3226 2753
rect 3282 2749 3286 2753
rect 3240 2740 3244 2747
rect 3298 2740 3302 2747
rect 3319 2744 3323 2748
rect 3336 2747 3340 2751
rect 3354 2749 3358 2753
rect 3414 2749 3418 2753
rect 3372 2740 3376 2747
rect 3430 2740 3434 2747
rect 3451 2744 3455 2748
rect 2001 2726 2005 2730
rect 2038 2724 2042 2728
rect 2058 2724 2062 2728
rect 2094 2724 2098 2728
rect 2133 2726 2137 2730
rect 2170 2724 2174 2728
rect 2190 2724 2194 2728
rect 2226 2724 2230 2728
rect 2265 2726 2269 2730
rect 2302 2724 2306 2728
rect 2322 2724 2326 2728
rect 2358 2724 2362 2728
rect 2397 2726 2401 2730
rect 2434 2724 2438 2728
rect 2454 2724 2458 2728
rect 2490 2724 2494 2728
rect 2946 2726 2950 2730
rect 2983 2724 2987 2728
rect 3003 2724 3007 2728
rect 3039 2724 3043 2728
rect 3078 2726 3082 2730
rect 3115 2724 3119 2728
rect 3135 2724 3139 2728
rect 3171 2724 3175 2728
rect 3210 2726 3214 2730
rect 3247 2724 3251 2728
rect 3267 2724 3271 2728
rect 3303 2724 3307 2728
rect 3342 2726 3346 2730
rect 3379 2724 3383 2728
rect 3399 2724 3403 2728
rect 3435 2724 3439 2728
rect 1643 2714 1647 2718
rect 1661 2716 1665 2720
rect 1721 2716 1725 2720
rect 1679 2707 1683 2714
rect 1737 2707 1741 2714
rect 1756 2711 1760 2715
rect 2588 2714 2592 2718
rect 2606 2716 2610 2720
rect 2666 2716 2670 2720
rect 2624 2707 2628 2714
rect 2682 2707 2686 2714
rect 2701 2711 2705 2715
rect 1649 2693 1653 2697
rect 1686 2691 1690 2695
rect 1706 2691 1710 2695
rect 1742 2691 1746 2695
rect 2017 2683 2021 2687
rect 2061 2683 2065 2687
rect 2088 2683 2092 2687
rect 2133 2683 2137 2687
rect 2206 2690 2210 2694
rect 1767 2670 1771 2674
rect 2171 2676 2175 2680
rect 1650 2661 1654 2665
rect 1997 2663 2001 2667
rect 2029 2664 2033 2668
rect 2048 2663 2052 2667
rect 2104 2664 2108 2668
rect 2120 2663 2124 2667
rect 2147 2663 2151 2667
rect 2287 2690 2291 2694
rect 2594 2693 2598 2697
rect 2198 2672 2202 2676
rect 2225 2668 2229 2672
rect 2252 2676 2256 2680
rect 2631 2691 2635 2695
rect 2651 2691 2655 2695
rect 2687 2691 2691 2695
rect 2279 2672 2283 2676
rect 2306 2668 2310 2672
rect 2962 2683 2966 2687
rect 3006 2683 3010 2687
rect 3033 2683 3037 2687
rect 3078 2683 3082 2687
rect 3151 2690 3155 2694
rect 2712 2670 2716 2674
rect 3116 2676 3120 2680
rect 2204 2654 2208 2658
rect 2595 2661 2599 2665
rect 2942 2663 2946 2667
rect 2285 2654 2289 2658
rect 2974 2664 2978 2668
rect 2993 2663 2997 2667
rect 3049 2664 3053 2668
rect 3065 2663 3069 2667
rect 3092 2663 3096 2667
rect 3232 2690 3236 2694
rect 3143 2672 3147 2676
rect 3170 2668 3174 2672
rect 3197 2676 3201 2680
rect 3224 2672 3228 2676
rect 3251 2668 3255 2672
rect 3149 2654 3153 2658
rect 3230 2654 3234 2658
rect 2014 2646 2018 2650
rect 2058 2645 2062 2649
rect 2083 2646 2088 2650
rect 2130 2645 2134 2649
rect 2959 2646 2963 2650
rect 3003 2645 3007 2649
rect 3028 2646 3033 2650
rect 3075 2645 3079 2649
rect 1649 2632 1653 2636
rect 1687 2632 1691 2636
rect 1707 2632 1711 2636
rect 1744 2632 1748 2636
rect 2594 2632 2598 2636
rect 2632 2632 2636 2636
rect 2652 2632 2656 2636
rect 2689 2632 2693 2636
rect 1637 2609 1641 2613
rect 1672 2614 1676 2618
rect 1656 2605 1660 2612
rect 1714 2605 1718 2612
rect 1732 2614 1736 2618
rect 2014 2616 2018 2620
rect 2058 2617 2062 2621
rect 1750 2612 1754 2616
rect 2083 2616 2088 2620
rect 2130 2617 2134 2621
rect 2206 2614 2210 2618
rect 2287 2614 2291 2618
rect 1997 2599 2001 2603
rect 1651 2589 1655 2593
rect 1687 2589 1691 2593
rect 1707 2589 1711 2593
rect 1744 2591 1748 2595
rect 2029 2598 2033 2602
rect 2048 2599 2052 2603
rect 2104 2598 2108 2602
rect 2120 2599 2124 2603
rect 2147 2599 2151 2603
rect 2195 2598 2201 2602
rect 2276 2598 2282 2602
rect 2582 2609 2586 2613
rect 2617 2614 2621 2618
rect 2601 2605 2605 2612
rect 2659 2605 2663 2612
rect 2677 2614 2681 2618
rect 2959 2616 2963 2620
rect 3003 2617 3007 2621
rect 2695 2612 2699 2616
rect 3028 2616 3033 2620
rect 3075 2617 3079 2621
rect 3151 2614 3155 2618
rect 3232 2614 3236 2618
rect 2942 2599 2946 2603
rect 2596 2589 2600 2593
rect 2632 2589 2636 2593
rect 2652 2589 2656 2593
rect 2689 2591 2693 2595
rect 2974 2598 2978 2602
rect 2993 2599 2997 2603
rect 3049 2598 3053 2602
rect 3065 2599 3069 2603
rect 3092 2599 3096 2603
rect 3140 2598 3146 2602
rect 3221 2598 3227 2602
rect 2017 2579 2021 2583
rect 2061 2579 2065 2583
rect 2088 2579 2092 2583
rect 2133 2579 2137 2583
rect 2204 2578 2208 2582
rect 2285 2578 2289 2582
rect 2962 2579 2966 2583
rect 3006 2579 3010 2583
rect 3033 2579 3037 2583
rect 3078 2579 3082 2583
rect 3149 2578 3153 2582
rect 3230 2578 3234 2582
rect 2206 2558 2210 2562
rect 2017 2551 2021 2555
rect 2061 2551 2065 2555
rect 2088 2551 2092 2555
rect 2133 2551 2137 2555
rect 2311 2558 2315 2562
rect 2198 2540 2202 2544
rect 1997 2531 2001 2535
rect 2029 2532 2033 2536
rect 2048 2531 2052 2535
rect 2104 2532 2108 2536
rect 2120 2531 2124 2535
rect 2147 2531 2151 2535
rect 2225 2536 2229 2540
rect 2276 2544 2280 2548
rect 3151 2558 3155 2562
rect 2303 2540 2307 2544
rect 2330 2536 2334 2540
rect 2962 2551 2966 2555
rect 3006 2551 3010 2555
rect 3033 2551 3037 2555
rect 3078 2551 3082 2555
rect 3256 2558 3260 2562
rect 3143 2540 3147 2544
rect 2942 2531 2946 2535
rect 2204 2522 2208 2526
rect 2309 2522 2313 2526
rect 2974 2532 2978 2536
rect 2993 2531 2997 2535
rect 3049 2532 3053 2536
rect 3065 2531 3069 2535
rect 3092 2531 3096 2535
rect 3170 2536 3174 2540
rect 3221 2544 3225 2548
rect 3248 2540 3252 2544
rect 3275 2536 3279 2540
rect 3149 2522 3153 2526
rect 3254 2522 3258 2526
rect 2014 2514 2018 2518
rect 2058 2513 2062 2517
rect 2083 2514 2088 2518
rect 2130 2513 2134 2517
rect 2959 2514 2963 2518
rect 3003 2513 3007 2517
rect 3028 2514 3033 2518
rect 3075 2513 3079 2517
rect 2014 2484 2018 2488
rect 2058 2485 2062 2489
rect 2083 2484 2088 2488
rect 2130 2485 2134 2489
rect 2206 2483 2210 2487
rect 2311 2483 2315 2487
rect 2959 2484 2963 2488
rect 3003 2485 3007 2489
rect 3028 2484 3033 2488
rect 3075 2485 3079 2489
rect 3151 2483 3155 2487
rect 3256 2483 3260 2487
rect 1997 2467 2001 2471
rect 2029 2466 2033 2470
rect 2048 2467 2052 2471
rect 2104 2466 2108 2470
rect 2120 2467 2124 2471
rect 2147 2467 2151 2471
rect 2195 2467 2201 2471
rect 2300 2467 2306 2471
rect 2942 2467 2946 2471
rect 2974 2466 2978 2470
rect 2993 2467 2997 2471
rect 3049 2466 3053 2470
rect 3065 2467 3069 2471
rect 3092 2467 3096 2471
rect 3140 2467 3146 2471
rect 3245 2467 3251 2471
rect 2017 2447 2021 2451
rect 2061 2447 2065 2451
rect 2088 2447 2092 2451
rect 2133 2447 2137 2451
rect 2204 2447 2208 2451
rect 2309 2447 2313 2451
rect 2962 2447 2966 2451
rect 3006 2447 3010 2451
rect 3033 2447 3037 2451
rect 3078 2447 3082 2451
rect 3149 2447 3153 2451
rect 3254 2447 3258 2451
rect 2206 2426 2210 2430
rect 2017 2419 2021 2423
rect 2061 2419 2065 2423
rect 2088 2419 2092 2423
rect 2133 2419 2137 2423
rect 2287 2426 2291 2430
rect 2198 2408 2202 2412
rect 1997 2399 2001 2403
rect 2029 2400 2033 2404
rect 2048 2399 2052 2403
rect 2104 2400 2108 2404
rect 2120 2399 2124 2403
rect 2147 2399 2151 2403
rect 2225 2404 2229 2408
rect 2252 2412 2256 2416
rect 2377 2426 2381 2430
rect 2279 2408 2283 2412
rect 2306 2404 2310 2408
rect 2342 2412 2346 2416
rect 3151 2426 3155 2430
rect 2369 2408 2373 2412
rect 2396 2404 2400 2408
rect 2962 2419 2966 2423
rect 3006 2419 3010 2423
rect 3033 2419 3037 2423
rect 3078 2419 3082 2423
rect 3232 2426 3236 2430
rect 3143 2408 3147 2412
rect 2942 2399 2946 2403
rect 2204 2390 2208 2394
rect 2285 2390 2289 2394
rect 2375 2390 2379 2394
rect 2974 2400 2978 2404
rect 2993 2399 2997 2403
rect 3049 2400 3053 2404
rect 3065 2399 3069 2403
rect 3092 2399 3096 2403
rect 3170 2404 3174 2408
rect 3197 2412 3201 2416
rect 3322 2426 3326 2430
rect 3224 2408 3228 2412
rect 3251 2404 3255 2408
rect 3287 2412 3291 2416
rect 3314 2408 3318 2412
rect 3341 2404 3345 2408
rect 3149 2390 3153 2394
rect 3230 2390 3234 2394
rect 3320 2390 3324 2394
rect 2014 2382 2018 2386
rect 2058 2381 2062 2385
rect 2083 2382 2088 2386
rect 2130 2381 2134 2385
rect 2959 2382 2963 2386
rect 3003 2381 3007 2385
rect 3028 2382 3033 2386
rect 3075 2381 3079 2385
rect 2014 2352 2018 2356
rect 2058 2353 2062 2357
rect 2083 2352 2088 2356
rect 2130 2353 2134 2357
rect 2959 2352 2963 2356
rect 3003 2353 3007 2357
rect 2206 2348 2210 2352
rect 2287 2348 2291 2352
rect 2377 2348 2381 2352
rect 3028 2352 3033 2356
rect 3075 2353 3079 2357
rect 3151 2348 3155 2352
rect 3232 2348 3236 2352
rect 3322 2348 3326 2352
rect 1997 2335 2001 2339
rect 2029 2334 2033 2338
rect 2048 2335 2052 2339
rect 2104 2334 2108 2338
rect 2120 2335 2124 2339
rect 2147 2335 2151 2339
rect 2195 2332 2201 2336
rect 2276 2332 2282 2336
rect 2366 2332 2372 2336
rect 2942 2335 2946 2339
rect 2974 2334 2978 2338
rect 2993 2335 2997 2339
rect 3049 2334 3053 2338
rect 3065 2335 3069 2339
rect 3092 2335 3096 2339
rect 3140 2332 3146 2336
rect 3221 2332 3227 2336
rect 3311 2332 3317 2336
rect 2017 2315 2021 2319
rect 2061 2315 2065 2319
rect 2088 2315 2092 2319
rect 2133 2315 2137 2319
rect 2204 2312 2208 2316
rect 2285 2312 2289 2316
rect 2375 2312 2379 2316
rect 2962 2315 2966 2319
rect 3006 2315 3010 2319
rect 3033 2315 3037 2319
rect 3078 2315 3082 2319
rect 3149 2312 3153 2316
rect 3230 2312 3234 2316
rect 3320 2312 3324 2316
rect 2206 2294 2210 2298
rect 2017 2287 2021 2291
rect 2061 2287 2065 2291
rect 2088 2287 2092 2291
rect 2133 2287 2137 2291
rect 3151 2294 3155 2298
rect 2198 2276 2202 2280
rect 1997 2267 2001 2271
rect 2029 2268 2033 2272
rect 2048 2267 2052 2271
rect 2104 2268 2108 2272
rect 2120 2267 2124 2271
rect 2147 2267 2151 2271
rect 2225 2272 2229 2276
rect 2962 2287 2966 2291
rect 3006 2287 3010 2291
rect 3033 2287 3037 2291
rect 3078 2287 3082 2291
rect 3143 2276 3147 2280
rect 2942 2267 2946 2271
rect 2204 2258 2208 2262
rect 2974 2268 2978 2272
rect 2993 2267 2997 2271
rect 3049 2268 3053 2272
rect 3065 2267 3069 2271
rect 3092 2267 3096 2271
rect 3170 2272 3174 2276
rect 3149 2258 3153 2262
rect 2014 2250 2018 2254
rect 2058 2249 2062 2253
rect 2083 2250 2088 2254
rect 2130 2249 2134 2253
rect 2959 2250 2963 2254
rect 3003 2249 3007 2253
rect 3028 2250 3033 2254
rect 3075 2249 3079 2253
rect 1517 2232 1521 2236
rect 1554 2232 1558 2236
rect 1574 2232 1578 2236
rect 1612 2232 1616 2236
rect 1649 2232 1653 2236
rect 1686 2232 1690 2236
rect 1706 2232 1710 2236
rect 1744 2232 1748 2236
rect 1781 2232 1785 2236
rect 1818 2232 1822 2236
rect 1838 2232 1842 2236
rect 1876 2232 1880 2236
rect 2462 2232 2466 2236
rect 2499 2232 2503 2236
rect 2519 2232 2523 2236
rect 2557 2232 2561 2236
rect 2594 2232 2598 2236
rect 2631 2232 2635 2236
rect 2651 2232 2655 2236
rect 2689 2232 2693 2236
rect 2726 2232 2730 2236
rect 2763 2232 2767 2236
rect 2783 2232 2787 2236
rect 2821 2232 2825 2236
rect 1511 2212 1515 2216
rect 1529 2214 1533 2218
rect 1589 2214 1593 2218
rect 1547 2205 1551 2212
rect 1605 2205 1609 2212
rect 1624 2209 1628 2213
rect 1642 2214 1646 2218
rect 1661 2214 1665 2218
rect 1721 2214 1725 2218
rect 1679 2205 1683 2212
rect 1737 2205 1741 2212
rect 1756 2209 1760 2213
rect 1774 2214 1778 2218
rect 1793 2214 1797 2218
rect 1853 2214 1857 2218
rect 1811 2205 1815 2212
rect 2014 2220 2018 2224
rect 2058 2221 2062 2225
rect 2083 2220 2088 2224
rect 2130 2221 2134 2225
rect 2275 2220 2279 2224
rect 2319 2221 2323 2225
rect 2344 2220 2349 2224
rect 2391 2221 2395 2225
rect 1869 2205 1873 2212
rect 1890 2209 1894 2213
rect 2206 2212 2210 2216
rect 2456 2212 2460 2216
rect 2474 2214 2478 2218
rect 1997 2203 2001 2207
rect 2029 2202 2033 2206
rect 2048 2203 2052 2207
rect 2104 2202 2108 2206
rect 2120 2203 2124 2207
rect 2147 2203 2151 2207
rect 1517 2191 1521 2195
rect 1554 2189 1558 2193
rect 1574 2189 1578 2193
rect 1610 2189 1614 2193
rect 1649 2191 1653 2195
rect 1686 2189 1690 2193
rect 1706 2189 1710 2193
rect 1742 2189 1746 2193
rect 1781 2191 1785 2195
rect 1818 2189 1822 2193
rect 1838 2189 1842 2193
rect 1874 2189 1878 2193
rect 2195 2196 2201 2200
rect 2233 2203 2237 2207
rect 2290 2202 2294 2206
rect 2309 2203 2313 2207
rect 2365 2202 2369 2206
rect 2381 2203 2385 2207
rect 2408 2203 2412 2207
rect 2534 2214 2538 2218
rect 2492 2205 2496 2212
rect 2550 2205 2554 2212
rect 2569 2209 2573 2213
rect 2587 2214 2591 2218
rect 2606 2214 2610 2218
rect 2666 2214 2670 2218
rect 2624 2205 2628 2212
rect 2682 2205 2686 2212
rect 2701 2209 2705 2213
rect 2719 2214 2723 2218
rect 2738 2214 2742 2218
rect 2798 2214 2802 2218
rect 2756 2205 2760 2212
rect 2959 2220 2963 2224
rect 3003 2221 3007 2225
rect 3028 2220 3033 2224
rect 3075 2221 3079 2225
rect 3220 2220 3224 2224
rect 3264 2221 3268 2225
rect 3289 2220 3294 2224
rect 3336 2221 3340 2225
rect 2814 2205 2818 2212
rect 2835 2209 2839 2213
rect 3151 2212 3155 2216
rect 2942 2203 2946 2207
rect 2974 2202 2978 2206
rect 2993 2203 2997 2207
rect 3049 2202 3053 2206
rect 3065 2203 3069 2207
rect 3092 2203 3096 2207
rect 2017 2183 2021 2187
rect 2061 2183 2065 2187
rect 2088 2183 2092 2187
rect 2133 2183 2137 2187
rect 2462 2191 2466 2195
rect 2204 2176 2208 2180
rect 1626 2161 1630 2165
rect 1650 2161 1654 2165
rect 2499 2189 2503 2193
rect 2519 2189 2523 2193
rect 2555 2189 2559 2193
rect 2594 2191 2598 2195
rect 2631 2189 2635 2193
rect 2651 2189 2655 2193
rect 2687 2189 2691 2193
rect 2726 2191 2730 2195
rect 2763 2189 2767 2193
rect 2783 2189 2787 2193
rect 2819 2189 2823 2193
rect 3140 2196 3146 2200
rect 3178 2203 3182 2207
rect 3235 2202 3239 2206
rect 3254 2203 3258 2207
rect 3310 2202 3314 2206
rect 3326 2203 3330 2207
rect 3353 2203 3357 2207
rect 2278 2183 2282 2187
rect 2322 2183 2326 2187
rect 2349 2183 2353 2187
rect 2394 2183 2398 2187
rect 2962 2183 2966 2187
rect 3006 2183 3010 2187
rect 3033 2183 3037 2187
rect 3078 2183 3082 2187
rect 3149 2176 3153 2180
rect 2571 2161 2575 2165
rect 2595 2161 2599 2165
rect 2417 2155 2421 2159
rect 2255 2148 2259 2152
rect 3223 2183 3227 2187
rect 3267 2183 3271 2187
rect 3294 2183 3298 2187
rect 3339 2183 3343 2187
rect 3362 2155 3366 2159
rect 3198 2148 3202 2152
rect 1646 2134 1650 2138
rect 2591 2134 2595 2138
rect 1661 2126 1665 2130
rect 2606 2126 2610 2130
rect 2300 2120 2304 2124
rect 2337 2120 2341 2124
rect 2357 2120 2361 2124
rect 2395 2120 2399 2124
rect 3245 2120 3249 2124
rect 3282 2120 3286 2124
rect 3302 2120 3306 2124
rect 3340 2120 3344 2124
rect 1626 2111 1630 2115
rect 1650 2111 1654 2115
rect 2571 2111 2575 2115
rect 2595 2111 2599 2115
rect 2294 2100 2298 2104
rect 2312 2102 2316 2106
rect 1517 2090 1521 2094
rect 1554 2090 1558 2094
rect 1574 2090 1578 2094
rect 1612 2090 1616 2094
rect 1649 2090 1653 2094
rect 1686 2090 1690 2094
rect 1706 2090 1710 2094
rect 1744 2090 1748 2094
rect 1781 2090 1785 2094
rect 1818 2090 1822 2094
rect 1838 2090 1842 2094
rect 1876 2090 1880 2094
rect 2372 2102 2376 2106
rect 2330 2093 2334 2100
rect 2388 2093 2392 2100
rect 2407 2097 2411 2101
rect 3239 2100 3243 2104
rect 3257 2102 3261 2106
rect 2462 2090 2466 2094
rect 2499 2090 2503 2094
rect 2519 2090 2523 2094
rect 2557 2090 2561 2094
rect 2594 2090 2598 2094
rect 2631 2090 2635 2094
rect 2651 2090 2655 2094
rect 2689 2090 2693 2094
rect 2726 2090 2730 2094
rect 2763 2090 2767 2094
rect 2783 2090 2787 2094
rect 2821 2090 2825 2094
rect 3317 2102 3321 2106
rect 3275 2093 3279 2100
rect 3333 2093 3337 2100
rect 3352 2097 3356 2101
rect 2300 2079 2304 2083
rect 1511 2070 1515 2074
rect 1529 2072 1533 2076
rect 1589 2072 1593 2076
rect 1547 2063 1551 2070
rect 1605 2063 1609 2070
rect 1624 2067 1628 2071
rect 1642 2072 1646 2076
rect 1661 2072 1665 2076
rect 1721 2072 1725 2076
rect 1679 2063 1683 2070
rect 1737 2063 1741 2070
rect 1756 2067 1760 2071
rect 1774 2072 1778 2076
rect 1793 2072 1797 2076
rect 1853 2072 1857 2076
rect 1811 2063 1815 2070
rect 2337 2077 2341 2081
rect 2357 2077 2361 2081
rect 2393 2077 2397 2081
rect 3245 2079 3249 2083
rect 1869 2063 1873 2070
rect 1890 2067 1894 2071
rect 2456 2070 2460 2074
rect 2474 2072 2478 2076
rect 2534 2072 2538 2076
rect 2492 2063 2496 2070
rect 2550 2063 2554 2070
rect 2569 2067 2573 2071
rect 2587 2072 2591 2076
rect 2606 2072 2610 2076
rect 2666 2072 2670 2076
rect 2624 2063 2628 2070
rect 2682 2063 2686 2070
rect 2701 2067 2705 2071
rect 2719 2072 2723 2076
rect 2738 2072 2742 2076
rect 2798 2072 2802 2076
rect 2756 2063 2760 2070
rect 3282 2077 3286 2081
rect 3302 2077 3306 2081
rect 3338 2077 3342 2081
rect 2814 2063 2818 2070
rect 2835 2067 2839 2071
rect 1517 2049 1521 2053
rect 1554 2047 1558 2051
rect 1574 2047 1578 2051
rect 1610 2047 1614 2051
rect 1649 2049 1653 2053
rect 1686 2047 1690 2051
rect 1706 2047 1710 2051
rect 1742 2047 1746 2051
rect 1781 2049 1785 2053
rect 1818 2047 1822 2051
rect 1838 2047 1842 2051
rect 1874 2047 1878 2051
rect 2462 2049 2466 2053
rect 2499 2047 2503 2051
rect 2519 2047 2523 2051
rect 2555 2047 2559 2051
rect 2594 2049 2598 2053
rect 2631 2047 2635 2051
rect 2651 2047 2655 2051
rect 2687 2047 2691 2051
rect 2726 2049 2730 2053
rect 2763 2047 2767 2051
rect 2783 2047 2787 2051
rect 2819 2047 2823 2051
rect 2300 2034 2304 2038
rect 2337 2034 2341 2038
rect 2357 2034 2361 2038
rect 2395 2034 2399 2038
rect 3245 2034 3249 2038
rect 3282 2034 3286 2038
rect 3302 2034 3306 2038
rect 3340 2034 3344 2038
rect 2294 2014 2298 2018
rect 2312 2016 2316 2020
rect 1517 2004 1521 2008
rect 1554 2004 1558 2008
rect 1574 2004 1578 2008
rect 1612 2004 1616 2008
rect 1649 2004 1653 2008
rect 1686 2004 1690 2008
rect 1706 2004 1710 2008
rect 1744 2004 1748 2008
rect 1781 2004 1785 2008
rect 1818 2004 1822 2008
rect 1838 2004 1842 2008
rect 1876 2004 1880 2008
rect 2372 2016 2376 2020
rect 2330 2007 2334 2014
rect 2388 2007 2392 2014
rect 2407 2011 2411 2015
rect 2429 2009 2433 2013
rect 3239 2014 3243 2018
rect 3257 2016 3261 2020
rect 2462 2004 2466 2008
rect 2499 2004 2503 2008
rect 2519 2004 2523 2008
rect 2557 2004 2561 2008
rect 2594 2004 2598 2008
rect 2631 2004 2635 2008
rect 2651 2004 2655 2008
rect 2689 2004 2693 2008
rect 2726 2004 2730 2008
rect 2763 2004 2767 2008
rect 2783 2004 2787 2008
rect 2821 2004 2825 2008
rect 3317 2016 3321 2020
rect 3275 2007 3279 2014
rect 3333 2007 3337 2014
rect 3352 2011 3356 2015
rect 3374 2009 3378 2013
rect 2300 1993 2304 1997
rect 1511 1984 1515 1988
rect 1529 1986 1533 1990
rect 1589 1986 1593 1990
rect 1547 1977 1551 1984
rect 1605 1977 1609 1984
rect 1624 1981 1628 1985
rect 1642 1986 1646 1990
rect 1661 1986 1665 1990
rect 1721 1986 1725 1990
rect 1679 1977 1683 1984
rect 1737 1977 1741 1984
rect 1756 1981 1760 1985
rect 1774 1986 1778 1990
rect 1793 1986 1797 1990
rect 1853 1986 1857 1990
rect 1811 1977 1815 1984
rect 2337 1991 2341 1995
rect 2357 1991 2361 1995
rect 2393 1991 2397 1995
rect 3245 1993 3249 1997
rect 1869 1977 1873 1984
rect 1890 1981 1894 1985
rect 2456 1984 2460 1988
rect 2474 1986 2478 1990
rect 2534 1986 2538 1990
rect 2492 1977 2496 1984
rect 2550 1977 2554 1984
rect 2569 1981 2573 1985
rect 2587 1986 2591 1990
rect 2606 1986 2610 1990
rect 2666 1986 2670 1990
rect 2624 1977 2628 1984
rect 2682 1977 2686 1984
rect 2701 1981 2705 1985
rect 2719 1986 2723 1990
rect 2738 1986 2742 1990
rect 2798 1986 2802 1990
rect 2756 1977 2760 1984
rect 3282 1991 3286 1995
rect 3302 1991 3306 1995
rect 3338 1991 3342 1995
rect 2814 1977 2818 1984
rect 2835 1981 2839 1985
rect 1517 1963 1521 1967
rect 1554 1961 1558 1965
rect 1574 1961 1578 1965
rect 1610 1961 1614 1965
rect 1649 1963 1653 1967
rect 1686 1961 1690 1965
rect 1706 1961 1710 1965
rect 1742 1961 1746 1965
rect 1781 1963 1785 1967
rect 1818 1961 1822 1965
rect 1838 1961 1842 1965
rect 1874 1961 1878 1965
rect 2462 1963 2466 1967
rect 2499 1961 2503 1965
rect 2519 1961 2523 1965
rect 2555 1961 2559 1965
rect 2594 1963 2598 1967
rect 2631 1961 2635 1965
rect 2651 1961 2655 1965
rect 2687 1961 2691 1965
rect 2726 1963 2730 1967
rect 2763 1961 2767 1965
rect 2783 1961 2787 1965
rect 2819 1961 2823 1965
rect 1743 1933 1747 1937
rect 1767 1933 1771 1937
rect 2688 1933 2692 1937
rect 2712 1933 2716 1937
rect 1763 1908 1767 1912
rect 2708 1908 2712 1912
rect 1778 1900 1782 1904
rect 2723 1900 2727 1904
rect 1743 1885 1747 1889
rect 1767 1885 1771 1889
rect 2688 1885 2692 1889
rect 2712 1885 2716 1889
rect 1517 1864 1521 1868
rect 1554 1864 1558 1868
rect 1574 1864 1578 1868
rect 1612 1864 1616 1868
rect 1649 1864 1653 1868
rect 1686 1864 1690 1868
rect 1706 1864 1710 1868
rect 1744 1864 1748 1868
rect 1781 1864 1785 1868
rect 1818 1864 1822 1868
rect 1838 1864 1842 1868
rect 1876 1864 1880 1868
rect 2462 1864 2466 1868
rect 2499 1864 2503 1868
rect 2519 1864 2523 1868
rect 2557 1864 2561 1868
rect 2594 1864 2598 1868
rect 2631 1864 2635 1868
rect 2651 1864 2655 1868
rect 2689 1864 2693 1868
rect 2726 1864 2730 1868
rect 2763 1864 2767 1868
rect 2783 1864 2787 1868
rect 2821 1864 2825 1868
rect 1511 1844 1515 1848
rect 1529 1846 1533 1850
rect 1589 1846 1593 1850
rect 1547 1837 1551 1844
rect 1605 1837 1609 1844
rect 1624 1841 1628 1845
rect 1642 1846 1646 1850
rect 1661 1846 1665 1850
rect 1721 1846 1725 1850
rect 1679 1837 1683 1844
rect 1737 1837 1741 1844
rect 1756 1841 1760 1845
rect 1774 1846 1778 1850
rect 1793 1846 1797 1850
rect 1853 1846 1857 1850
rect 1811 1837 1815 1844
rect 1869 1837 1873 1844
rect 1890 1841 1894 1845
rect 2456 1844 2460 1848
rect 2474 1846 2478 1850
rect 2534 1846 2538 1850
rect 2492 1837 2496 1844
rect 2550 1837 2554 1844
rect 2569 1841 2573 1845
rect 2587 1846 2591 1850
rect 2606 1846 2610 1850
rect 2666 1846 2670 1850
rect 2624 1837 2628 1844
rect 2682 1837 2686 1844
rect 2701 1841 2705 1845
rect 2719 1846 2723 1850
rect 2738 1846 2742 1850
rect 2798 1846 2802 1850
rect 2756 1837 2760 1844
rect 2814 1837 2818 1844
rect 2835 1841 2839 1845
rect 1517 1823 1521 1827
rect 1554 1821 1558 1825
rect 1574 1821 1578 1825
rect 1610 1821 1614 1825
rect 1649 1823 1653 1827
rect 1686 1821 1690 1825
rect 1706 1821 1710 1825
rect 1742 1821 1746 1825
rect 1781 1823 1785 1827
rect 1818 1821 1822 1825
rect 1838 1821 1842 1825
rect 1874 1821 1878 1825
rect 2462 1823 2466 1827
rect 2499 1821 2503 1825
rect 2519 1821 2523 1825
rect 2555 1821 2559 1825
rect 2594 1823 2598 1827
rect 2631 1821 2635 1825
rect 2651 1821 2655 1825
rect 2687 1821 2691 1825
rect 2726 1823 2730 1827
rect 2763 1821 2767 1825
rect 2783 1821 2787 1825
rect 2819 1821 2823 1825
<< metal1 >>
rect 1376 4845 1460 4930
rect 1679 4820 1757 4909
rect 1986 4825 2064 4914
rect 2303 4825 2381 4914
rect 2614 4827 2692 4916
rect 2918 4817 2996 4906
rect 3232 4825 3310 4914
rect 3522 4810 3634 4924
rect 1718 4300 1731 4326
rect 2027 4304 2040 4326
rect 2336 4304 2349 4354
rect 2645 4316 2658 4338
rect 2954 4303 2967 4338
rect 3263 4314 3276 4338
rect 2695 4298 2967 4303
rect 2994 4299 3279 4314
rect 3548 4289 3604 4336
rect 2958 4284 3604 4289
rect 2693 4280 2713 4284
rect 2717 4280 2767 4284
rect 2771 4280 2910 4284
rect 2914 4280 2962 4284
rect 2696 4276 2699 4280
rect 2705 4263 2708 4268
rect 2720 4270 2723 4280
rect 2750 4276 2753 4280
rect 2689 4259 2690 4262
rect 2694 4259 2697 4262
rect 2736 4259 2739 4262
rect 2705 4254 2708 4259
rect 2713 4255 2724 4258
rect 2736 4256 2744 4259
rect 2736 4250 2739 4256
rect 2748 4251 2751 4254
rect 2759 4254 2762 4268
rect 2870 4273 2873 4280
rect 2923 4273 2926 4280
rect 2759 4251 2771 4254
rect 2696 4204 2699 4250
rect 2759 4246 2762 4251
rect 2720 4204 2723 4246
rect 2750 4204 2753 4242
rect 2768 4236 2771 4251
rect 3002 4278 3126 4279
rect 3548 4278 3604 4284
rect 3002 4264 3605 4278
rect 3027 4263 3605 4264
rect 3881 4259 3894 4318
rect 3010 4246 3894 4259
rect 2768 4231 2885 4236
rect 2903 4235 2906 4243
rect 2956 4235 2959 4243
rect 2903 4231 2923 4235
rect 2927 4231 2938 4235
rect 2903 4223 2906 4231
rect 2956 4223 2959 4231
rect 2870 4204 2873 4211
rect 2923 4204 2926 4211
rect 2693 4200 2713 4204
rect 2717 4200 2767 4204
rect 2771 4200 2910 4204
rect 2914 4200 2990 4204
rect 2720 4190 2723 4200
rect 2660 4178 2721 4181
rect 2736 4180 2739 4186
rect 2736 4177 2744 4180
rect 2736 4174 2739 4177
rect 2720 4154 2723 4166
rect 2671 4150 2689 4154
rect 2693 4150 2713 4154
rect 2717 4150 2767 4154
rect 2771 4150 2816 4154
rect 2820 4150 2998 4154
rect 2674 4146 2677 4150
rect 2696 4146 2699 4150
rect 2683 4133 2686 4138
rect 2705 4133 2708 4138
rect 2720 4140 2723 4150
rect 2750 4146 2753 4150
rect 2667 4129 2668 4132
rect 2672 4129 2675 4132
rect 2687 4129 2690 4133
rect 2694 4129 2697 4132
rect 2736 4129 2739 4132
rect 2683 4124 2686 4129
rect 2705 4124 2708 4129
rect 2713 4125 2724 4128
rect 2736 4126 2744 4129
rect 2736 4120 2739 4126
rect 2748 4121 2751 4124
rect 2759 4124 2762 4138
rect 2776 4143 2779 4150
rect 2829 4143 2832 4150
rect 2759 4121 2771 4124
rect 2674 4074 2677 4120
rect 2696 4074 2699 4120
rect 2759 4116 2762 4121
rect 2720 4074 2723 4116
rect 2750 4074 2753 4112
rect 2768 4106 2771 4121
rect 2768 4101 2791 4106
rect 2809 4105 2812 4113
rect 2862 4106 2865 4113
rect 2809 4101 2818 4105
rect 2822 4101 2844 4105
rect 2809 4093 2812 4101
rect 2862 4093 2865 4102
rect 2776 4074 2779 4081
rect 2829 4074 2832 4081
rect 2671 4070 2689 4074
rect 2693 4070 2713 4074
rect 2717 4070 2767 4074
rect 2771 4070 2816 4074
rect 2820 4070 2990 4074
rect 2720 4060 2723 4070
rect 2662 4048 2721 4051
rect 2736 4050 2739 4056
rect 2736 4047 2744 4050
rect 2736 4044 2739 4047
rect 2720 4024 2723 4036
rect 2689 4020 2713 4024
rect 2717 4020 2998 4024
rect 2867 3994 2923 3998
rect 2879 3987 2930 3991
rect 1901 3962 2027 3966
rect 1991 3951 2336 3955
rect 1970 3943 2897 3947
rect 1958 3935 2885 3939
rect 1946 3928 2873 3932
rect 1934 3921 2861 3925
rect 1922 3913 2849 3917
rect 2855 3913 2990 3917
rect 2832 3909 2837 3910
rect 1910 3906 2837 3909
rect 2843 3906 2998 3910
rect 1910 3905 2838 3906
rect 1982 3898 2921 3902
rect 2927 3898 3006 3902
rect 2903 3836 2909 3840
rect 2891 3828 2897 3832
rect 2879 3820 2885 3824
rect 1620 3815 1897 3819
rect 2867 3812 2873 3816
rect 1642 3807 1987 3811
rect 2855 3804 2861 3808
rect 2843 3796 2849 3800
rect 1970 3763 1997 3767
rect 2001 3763 2033 3767
rect 2037 3763 2100 3767
rect 2104 3763 2129 3767
rect 2133 3763 2165 3767
rect 2169 3763 2232 3767
rect 2236 3763 2261 3767
rect 2265 3763 2297 3767
rect 2301 3763 2364 3767
rect 2368 3763 2393 3767
rect 2397 3763 2429 3767
rect 2433 3763 2496 3767
rect 2500 3763 2516 3767
rect 2915 3763 2942 3767
rect 2946 3763 2978 3767
rect 2982 3763 3045 3767
rect 3049 3763 3074 3767
rect 3078 3763 3110 3767
rect 3114 3763 3177 3767
rect 3181 3763 3206 3767
rect 3210 3763 3242 3767
rect 3246 3763 3309 3767
rect 3313 3763 3338 3767
rect 3342 3763 3374 3767
rect 3378 3763 3441 3767
rect 3445 3763 3461 3767
rect 1910 3756 2021 3760
rect 2025 3756 2049 3760
rect 2053 3756 2079 3760
rect 2083 3756 2116 3760
rect 2120 3756 2153 3760
rect 2157 3756 2181 3760
rect 2185 3756 2211 3760
rect 2215 3756 2248 3760
rect 2252 3756 2285 3760
rect 2289 3756 2313 3760
rect 2317 3756 2343 3760
rect 2347 3756 2380 3760
rect 2384 3756 2417 3760
rect 2421 3756 2445 3760
rect 2449 3756 2475 3760
rect 2479 3756 2512 3760
rect 2855 3756 2966 3760
rect 2970 3756 2994 3760
rect 2998 3756 3024 3760
rect 3028 3756 3061 3760
rect 3065 3756 3098 3760
rect 3102 3756 3126 3760
rect 3130 3756 3156 3760
rect 3160 3756 3193 3760
rect 3197 3756 3230 3760
rect 3234 3756 3258 3760
rect 3262 3756 3288 3760
rect 3292 3756 3325 3760
rect 3329 3756 3362 3760
rect 3366 3756 3390 3760
rect 3394 3756 3420 3760
rect 3424 3756 3457 3760
rect 1991 3746 1994 3756
rect 2012 3746 2015 3756
rect 2028 3746 2031 3756
rect 2042 3749 2047 3753
rect 2051 3749 2058 3753
rect 2070 3746 2073 3756
rect 2086 3746 2089 3756
rect 2107 3746 2110 3756
rect 2123 3746 2126 3756
rect 2144 3746 2147 3756
rect 2160 3746 2163 3756
rect 2174 3749 2179 3753
rect 2183 3749 2190 3753
rect 2202 3746 2205 3756
rect 2218 3746 2221 3756
rect 2239 3746 2242 3756
rect 2255 3746 2258 3756
rect 2276 3746 2279 3756
rect 2292 3746 2295 3756
rect 2306 3749 2311 3753
rect 2315 3749 2322 3753
rect 2334 3746 2337 3756
rect 2350 3746 2353 3756
rect 2371 3746 2374 3756
rect 2387 3746 2390 3756
rect 2408 3746 2411 3756
rect 2424 3746 2427 3756
rect 2438 3749 2443 3753
rect 2447 3749 2454 3753
rect 2466 3746 2469 3756
rect 2482 3746 2485 3756
rect 2503 3746 2506 3756
rect 2936 3746 2939 3756
rect 2957 3746 2960 3756
rect 2973 3746 2976 3756
rect 2987 3749 2992 3753
rect 2996 3749 3003 3753
rect 3015 3746 3018 3756
rect 3031 3746 3034 3756
rect 3052 3746 3055 3756
rect 3068 3746 3071 3756
rect 3089 3746 3092 3756
rect 3105 3746 3108 3756
rect 3119 3749 3124 3753
rect 3128 3749 3135 3753
rect 3147 3746 3150 3756
rect 3163 3746 3166 3756
rect 3184 3746 3187 3756
rect 3200 3746 3203 3756
rect 3221 3746 3224 3756
rect 3237 3746 3240 3756
rect 3251 3749 3256 3753
rect 3260 3749 3267 3753
rect 3279 3746 3282 3756
rect 3295 3746 3298 3756
rect 3316 3746 3319 3756
rect 3332 3746 3335 3756
rect 3353 3746 3356 3756
rect 3369 3746 3372 3756
rect 3383 3749 3388 3753
rect 3392 3749 3399 3753
rect 3411 3746 3414 3756
rect 3427 3746 3430 3756
rect 3448 3746 3451 3756
rect 1636 3730 1645 3734
rect 1649 3730 1681 3734
rect 1685 3730 1748 3734
rect 1752 3730 1964 3734
rect 2008 3732 2013 3735
rect 2017 3732 2041 3735
rect 2066 3732 2073 3735
rect 2077 3732 2099 3735
rect 1636 3723 1669 3727
rect 1673 3723 1697 3727
rect 1701 3723 1727 3727
rect 1731 3723 1764 3727
rect 1768 3723 1904 3727
rect 1639 3713 1642 3723
rect 1660 3713 1663 3723
rect 1676 3713 1679 3723
rect 1690 3716 1695 3720
rect 1699 3716 1706 3720
rect 1718 3713 1721 3723
rect 1734 3713 1737 3723
rect 1755 3713 1758 3723
rect 2024 3722 2031 3725
rect 2035 3726 2054 3729
rect 2054 3719 2057 3725
rect 2082 3722 2089 3725
rect 2093 3726 2110 3729
rect 2140 3732 2145 3735
rect 2149 3732 2173 3735
rect 2198 3732 2205 3735
rect 2209 3732 2231 3735
rect 2156 3722 2163 3725
rect 2167 3726 2186 3729
rect 2186 3719 2189 3725
rect 2214 3722 2221 3725
rect 2225 3726 2242 3729
rect 2272 3732 2277 3735
rect 2281 3732 2305 3735
rect 2330 3732 2337 3735
rect 2341 3732 2363 3735
rect 2288 3722 2295 3725
rect 2299 3726 2318 3729
rect 2318 3719 2321 3725
rect 2346 3722 2353 3725
rect 2357 3726 2374 3729
rect 2404 3732 2409 3735
rect 2413 3732 2437 3735
rect 2462 3732 2469 3735
rect 2473 3732 2495 3735
rect 2581 3730 2590 3734
rect 2594 3730 2626 3734
rect 2630 3730 2693 3734
rect 2697 3730 2909 3734
rect 2420 3722 2427 3725
rect 2431 3726 2450 3729
rect 1634 3696 1643 3700
rect 1656 3699 1661 3702
rect 1665 3699 1689 3702
rect 1714 3699 1721 3702
rect 1725 3699 1747 3702
rect 1991 3703 1994 3715
rect 2012 3703 2015 3715
rect 2028 3703 2031 3715
rect 2042 3706 2054 3709
rect 2070 3703 2073 3715
rect 2086 3703 2089 3715
rect 2107 3703 2110 3715
rect 2123 3703 2126 3715
rect 2144 3703 2147 3715
rect 2160 3703 2163 3715
rect 2174 3706 2186 3709
rect 2202 3703 2205 3715
rect 2218 3703 2221 3715
rect 2239 3703 2242 3715
rect 2255 3703 2258 3715
rect 2276 3703 2279 3715
rect 2292 3703 2295 3715
rect 2306 3706 2318 3709
rect 2334 3703 2337 3715
rect 2350 3703 2353 3715
rect 2371 3703 2374 3715
rect 2450 3719 2453 3725
rect 2478 3722 2485 3725
rect 2489 3726 2506 3729
rect 2953 3732 2958 3735
rect 2962 3732 2986 3735
rect 3011 3732 3018 3735
rect 3022 3732 3044 3735
rect 2581 3723 2614 3727
rect 2618 3723 2642 3727
rect 2646 3723 2672 3727
rect 2676 3723 2709 3727
rect 2713 3723 2849 3727
rect 2387 3703 2390 3715
rect 2408 3703 2411 3715
rect 2424 3703 2427 3715
rect 2438 3706 2450 3709
rect 2466 3703 2469 3715
rect 2482 3703 2485 3715
rect 2503 3703 2506 3715
rect 2584 3713 2587 3723
rect 2605 3713 2608 3723
rect 2621 3713 2624 3723
rect 2635 3716 2640 3720
rect 2644 3716 2651 3720
rect 2663 3713 2666 3723
rect 2679 3713 2682 3723
rect 2700 3713 2703 3723
rect 2969 3722 2976 3725
rect 2980 3726 2999 3729
rect 2999 3719 3002 3725
rect 3027 3722 3034 3725
rect 3038 3726 3055 3729
rect 3085 3732 3090 3735
rect 3094 3732 3118 3735
rect 3143 3732 3150 3735
rect 3154 3732 3176 3735
rect 3101 3722 3108 3725
rect 3112 3726 3131 3729
rect 3131 3719 3134 3725
rect 3159 3722 3166 3725
rect 3170 3726 3187 3729
rect 3217 3732 3222 3735
rect 3226 3732 3250 3735
rect 3275 3732 3282 3735
rect 3286 3732 3308 3735
rect 3233 3722 3240 3725
rect 3244 3726 3263 3729
rect 3263 3719 3266 3725
rect 3291 3722 3298 3725
rect 3302 3726 3319 3729
rect 3349 3732 3354 3735
rect 3358 3732 3382 3735
rect 3407 3732 3414 3735
rect 3418 3732 3440 3735
rect 3365 3722 3372 3725
rect 3376 3726 3395 3729
rect 1922 3699 2021 3703
rect 2025 3699 2049 3703
rect 2053 3699 2079 3703
rect 2083 3699 2153 3703
rect 2157 3699 2181 3703
rect 2185 3699 2211 3703
rect 2215 3699 2285 3703
rect 2289 3699 2313 3703
rect 2317 3699 2343 3703
rect 2347 3699 2417 3703
rect 2421 3699 2445 3703
rect 2449 3699 2475 3703
rect 2479 3699 2516 3703
rect 1672 3689 1679 3692
rect 1683 3693 1702 3696
rect 1702 3686 1705 3692
rect 1730 3689 1737 3692
rect 1741 3693 1756 3696
rect 2579 3696 2588 3700
rect 2601 3699 2606 3702
rect 2610 3699 2634 3702
rect 2659 3699 2666 3702
rect 2670 3699 2692 3702
rect 2936 3703 2939 3715
rect 2957 3703 2960 3715
rect 2973 3703 2976 3715
rect 2987 3706 2999 3709
rect 3015 3703 3018 3715
rect 3031 3703 3034 3715
rect 3052 3703 3055 3715
rect 3068 3703 3071 3715
rect 3089 3703 3092 3715
rect 3105 3703 3108 3715
rect 3119 3706 3131 3709
rect 3147 3703 3150 3715
rect 3163 3703 3166 3715
rect 3184 3703 3187 3715
rect 3200 3703 3203 3715
rect 3221 3703 3224 3715
rect 3237 3703 3240 3715
rect 3251 3706 3263 3709
rect 3279 3703 3282 3715
rect 3295 3703 3298 3715
rect 3316 3703 3319 3715
rect 3395 3719 3398 3725
rect 3423 3722 3430 3725
rect 3434 3726 3451 3729
rect 3332 3703 3335 3715
rect 3353 3703 3356 3715
rect 3369 3703 3372 3715
rect 3383 3706 3395 3709
rect 3411 3703 3414 3715
rect 3427 3703 3430 3715
rect 3448 3703 3451 3715
rect 2867 3699 2966 3703
rect 2970 3699 2994 3703
rect 2998 3699 3024 3703
rect 3028 3699 3098 3703
rect 3102 3699 3126 3703
rect 3130 3699 3156 3703
rect 3160 3699 3230 3703
rect 3234 3699 3258 3703
rect 3262 3699 3288 3703
rect 3292 3699 3362 3703
rect 3366 3699 3390 3703
rect 3394 3699 3420 3703
rect 3424 3699 3461 3703
rect 1958 3692 1997 3696
rect 2001 3692 2048 3696
rect 2052 3692 2098 3696
rect 2102 3692 2129 3696
rect 2133 3692 2180 3696
rect 2184 3692 2230 3696
rect 2234 3692 2261 3696
rect 2265 3692 2312 3696
rect 2316 3692 2362 3696
rect 2366 3692 2393 3696
rect 2397 3692 2444 3696
rect 2448 3692 2494 3696
rect 2498 3692 2516 3696
rect 2617 3689 2624 3692
rect 2628 3693 2647 3696
rect 1639 3670 1642 3682
rect 1660 3670 1663 3682
rect 1676 3670 1679 3682
rect 1690 3673 1702 3676
rect 1718 3670 1721 3682
rect 1734 3670 1737 3682
rect 1755 3670 1758 3682
rect 1910 3679 1995 3683
rect 1999 3679 2011 3683
rect 2015 3679 2029 3683
rect 2033 3679 2040 3683
rect 2044 3679 2046 3683
rect 2050 3679 2065 3683
rect 2069 3679 2102 3683
rect 2106 3679 2107 3683
rect 2111 3679 2119 3683
rect 2123 3679 2147 3683
rect 2151 3679 2163 3683
rect 2167 3679 2187 3683
rect 2191 3679 2241 3683
rect 2245 3679 2268 3683
rect 2272 3679 2322 3683
rect 2326 3679 2345 3683
rect 2647 3686 2650 3692
rect 2675 3689 2682 3692
rect 2686 3693 2701 3696
rect 2903 3692 2942 3696
rect 2946 3692 2993 3696
rect 2997 3692 3043 3696
rect 3047 3692 3074 3696
rect 3078 3692 3125 3696
rect 3129 3692 3175 3696
rect 3179 3692 3206 3696
rect 3210 3692 3257 3696
rect 3261 3692 3307 3696
rect 3311 3692 3338 3696
rect 3342 3692 3389 3696
rect 3393 3692 3439 3696
rect 3443 3692 3461 3696
rect 1946 3672 2022 3676
rect 2026 3672 2053 3676
rect 2057 3672 2075 3676
rect 2079 3672 2140 3676
rect 2144 3672 2158 3676
rect 2170 3675 2173 3679
rect 1636 3666 1669 3670
rect 1673 3666 1697 3670
rect 1701 3666 1727 3670
rect 1731 3666 1916 3670
rect 1636 3659 1645 3663
rect 1649 3659 1696 3663
rect 1700 3659 1746 3663
rect 1750 3659 1952 3663
rect 2065 3665 2068 3669
rect 2092 3665 2093 3669
rect 2137 3665 2139 3669
rect 2179 3662 2182 3667
rect 2194 3669 2197 3679
rect 2224 3675 2227 3679
rect 2251 3675 2254 3679
rect 1634 3643 1650 3647
rect 1759 3645 1763 3649
rect 1775 3645 1779 3649
rect 1783 3645 1997 3649
rect 2005 3648 2008 3654
rect 2012 3648 2015 3654
rect 2005 3645 2015 3648
rect 2005 3640 2008 3645
rect 1642 3636 1646 3640
rect 1658 3636 1779 3640
rect 2012 3640 2015 3645
rect 2021 3650 2024 3654
rect 2021 3646 2023 3650
rect 2027 3646 2029 3650
rect 2037 3649 2040 3654
rect 2065 3651 2068 3654
rect 2037 3647 2048 3649
rect 2021 3640 2024 3646
rect 2037 3645 2043 3647
rect 2037 3640 2040 3645
rect 2047 3645 2048 3647
rect 2066 3647 2068 3651
rect 2065 3640 2068 3647
rect 2168 3658 2171 3661
rect 2210 3658 2213 3661
rect 2081 3650 2084 3654
rect 2091 3650 2094 3654
rect 2091 3646 2100 3650
rect 2112 3649 2115 3654
rect 2137 3650 2140 3654
rect 2081 3640 2084 3646
rect 2091 3640 2094 3646
rect 2112 3645 2113 3649
rect 2117 3645 2120 3648
rect 2139 3646 2140 3650
rect 2155 3649 2158 3654
rect 2179 3653 2182 3658
rect 2187 3654 2198 3657
rect 2210 3655 2218 3658
rect 2112 3640 2115 3645
rect 2137 3640 2140 3646
rect 2155 3640 2158 3645
rect 1629 3628 1645 3632
rect 1649 3628 1712 3632
rect 1716 3628 1748 3632
rect 1752 3628 1964 3632
rect 2057 3627 2058 3631
rect 2082 3628 2083 3632
rect 2129 3627 2130 3631
rect 1633 3621 1666 3625
rect 1670 3621 1696 3625
rect 1700 3621 1724 3625
rect 1728 3621 1904 3625
rect 1639 3611 1642 3621
rect 1660 3611 1663 3621
rect 1676 3611 1679 3621
rect 1691 3614 1698 3618
rect 1702 3614 1707 3618
rect 1718 3611 1721 3621
rect 1734 3611 1737 3621
rect 1755 3611 1758 3621
rect 1934 3620 2010 3624
rect 2014 3620 2069 3624
rect 2073 3620 2094 3624
rect 2098 3620 2125 3624
rect 2129 3620 2158 3624
rect 2170 3617 2173 3649
rect 2187 3648 2190 3654
rect 2210 3649 2213 3655
rect 2222 3650 2225 3653
rect 2233 3653 2236 3667
rect 2260 3662 2263 3667
rect 2275 3669 2278 3679
rect 2305 3675 2308 3679
rect 2244 3658 2245 3661
rect 2249 3658 2252 3661
rect 2584 3670 2587 3682
rect 2605 3670 2608 3682
rect 2621 3670 2624 3682
rect 2635 3673 2647 3676
rect 2663 3670 2666 3682
rect 2679 3670 2682 3682
rect 2700 3670 2703 3682
rect 2855 3679 2940 3683
rect 2944 3679 2956 3683
rect 2960 3679 2974 3683
rect 2978 3679 2985 3683
rect 2989 3679 2991 3683
rect 2995 3679 3010 3683
rect 3014 3679 3047 3683
rect 3051 3679 3052 3683
rect 3056 3679 3064 3683
rect 3068 3679 3092 3683
rect 3096 3679 3108 3683
rect 3112 3679 3132 3683
rect 3136 3679 3186 3683
rect 3190 3679 3213 3683
rect 3217 3679 3267 3683
rect 3271 3679 3290 3683
rect 2891 3672 2967 3676
rect 2971 3672 2998 3676
rect 3002 3672 3020 3676
rect 3024 3672 3085 3676
rect 3089 3672 3103 3676
rect 3115 3675 3118 3679
rect 2291 3658 2294 3661
rect 2233 3650 2241 3653
rect 2260 3653 2263 3658
rect 2233 3645 2236 3650
rect 2241 3646 2245 3650
rect 2268 3654 2279 3657
rect 2291 3655 2299 3658
rect 2185 3639 2190 3644
rect 2194 3617 2197 3645
rect 2224 3617 2227 3641
rect 2251 3617 2254 3649
rect 2268 3648 2271 3654
rect 2291 3649 2294 3655
rect 2303 3650 2306 3653
rect 2314 3653 2317 3667
rect 2581 3666 2614 3670
rect 2618 3666 2642 3670
rect 2646 3666 2672 3670
rect 2676 3666 2861 3670
rect 2581 3659 2590 3663
rect 2594 3659 2641 3663
rect 2645 3659 2691 3663
rect 2695 3659 2897 3663
rect 3010 3665 3013 3669
rect 3037 3665 3038 3669
rect 3082 3665 3084 3669
rect 3124 3662 3127 3667
rect 3139 3669 3142 3679
rect 3169 3675 3172 3679
rect 3196 3675 3199 3679
rect 2314 3650 2326 3653
rect 2314 3645 2317 3650
rect 2266 3639 2271 3644
rect 2275 3617 2278 3645
rect 2579 3643 2595 3647
rect 2704 3645 2708 3649
rect 2720 3645 2724 3649
rect 2728 3645 2933 3649
rect 2937 3645 2942 3649
rect 2950 3648 2953 3654
rect 2957 3648 2960 3654
rect 2950 3645 2960 3648
rect 2305 3617 2308 3641
rect 2950 3640 2953 3645
rect 2587 3636 2591 3640
rect 2603 3636 2724 3640
rect 2957 3640 2960 3645
rect 2966 3650 2969 3654
rect 2966 3646 2968 3650
rect 2972 3646 2974 3650
rect 2982 3649 2985 3654
rect 3010 3651 3013 3654
rect 2982 3647 2993 3649
rect 2966 3640 2969 3646
rect 2982 3645 2988 3647
rect 2982 3640 2985 3645
rect 2992 3645 2993 3647
rect 3011 3647 3013 3651
rect 3010 3640 3013 3647
rect 3113 3658 3116 3661
rect 3155 3658 3158 3661
rect 3026 3650 3029 3654
rect 3036 3650 3039 3654
rect 3036 3646 3045 3650
rect 3057 3649 3060 3654
rect 3082 3650 3085 3654
rect 3026 3640 3029 3646
rect 3036 3640 3039 3646
rect 3057 3645 3058 3649
rect 3062 3645 3065 3648
rect 3084 3646 3085 3650
rect 3100 3649 3103 3654
rect 3124 3653 3127 3658
rect 3132 3654 3143 3657
rect 3155 3655 3163 3658
rect 3057 3640 3060 3645
rect 3082 3640 3085 3646
rect 3100 3640 3103 3645
rect 2574 3628 2590 3632
rect 2594 3628 2657 3632
rect 2661 3628 2693 3632
rect 2697 3628 2909 3632
rect 3002 3627 3003 3631
rect 3027 3628 3028 3632
rect 3074 3627 3075 3631
rect 2578 3621 2611 3625
rect 2615 3621 2641 3625
rect 2645 3621 2669 3625
rect 2673 3621 2849 3625
rect 1922 3613 1996 3617
rect 2000 3613 2002 3617
rect 2006 3613 2010 3617
rect 2014 3613 2028 3617
rect 2032 3613 2037 3617
rect 2041 3613 2046 3617
rect 2050 3613 2069 3617
rect 2073 3613 2103 3617
rect 2107 3613 2118 3617
rect 2122 3613 2146 3617
rect 2150 3613 2163 3617
rect 2167 3613 2187 3617
rect 2191 3613 2241 3617
rect 2248 3613 2268 3617
rect 2272 3613 2322 3617
rect 1650 3597 1672 3600
rect 1676 3597 1683 3600
rect 1934 3606 2010 3610
rect 2014 3606 2069 3610
rect 2073 3606 2094 3610
rect 2098 3606 2125 3610
rect 2129 3606 2158 3610
rect 1708 3597 1732 3600
rect 1736 3597 1741 3600
rect 2057 3599 2058 3603
rect 2082 3598 2083 3602
rect 2129 3599 2130 3603
rect 1754 3594 1763 3598
rect 1641 3591 1656 3594
rect 1695 3591 1714 3594
rect 1660 3587 1667 3590
rect 1692 3584 1695 3590
rect 1718 3587 1725 3590
rect 2005 3585 2008 3590
rect 2012 3585 2015 3590
rect 1995 3582 1997 3585
rect 2005 3582 2015 3585
rect 1639 3568 1642 3580
rect 1660 3568 1663 3580
rect 1676 3568 1679 3580
rect 1695 3571 1707 3574
rect 1718 3568 1721 3580
rect 1734 3568 1737 3580
rect 1755 3568 1758 3580
rect 2005 3576 2008 3582
rect 2012 3576 2015 3582
rect 2021 3584 2024 3590
rect 2037 3585 2040 3590
rect 2021 3580 2023 3584
rect 2027 3580 2029 3584
rect 2037 3583 2043 3585
rect 2047 3583 2048 3585
rect 2037 3581 2048 3583
rect 2065 3583 2068 3590
rect 2021 3576 2024 3580
rect 2037 3576 2040 3581
rect 2066 3579 2068 3583
rect 2065 3576 2068 3579
rect 2081 3584 2084 3590
rect 2091 3584 2094 3590
rect 2112 3585 2115 3590
rect 2091 3580 2100 3584
rect 2112 3581 2113 3585
rect 2117 3582 2120 3585
rect 2137 3584 2140 3590
rect 2155 3585 2158 3590
rect 2194 3593 2197 3613
rect 2275 3593 2278 3613
rect 2584 3611 2587 3621
rect 2605 3611 2608 3621
rect 2621 3611 2624 3621
rect 2636 3614 2643 3618
rect 2647 3614 2652 3618
rect 2663 3611 2666 3621
rect 2679 3611 2682 3621
rect 2700 3611 2703 3621
rect 2879 3620 2955 3624
rect 2959 3620 3014 3624
rect 3018 3620 3039 3624
rect 3043 3620 3070 3624
rect 3074 3620 3103 3624
rect 3115 3617 3118 3649
rect 3132 3648 3135 3654
rect 3155 3649 3158 3655
rect 3167 3650 3170 3653
rect 3178 3653 3181 3667
rect 3205 3662 3208 3667
rect 3220 3669 3223 3679
rect 3250 3675 3253 3679
rect 3189 3658 3190 3661
rect 3194 3658 3197 3661
rect 3236 3658 3239 3661
rect 3178 3650 3186 3653
rect 3205 3653 3208 3658
rect 3178 3645 3181 3650
rect 3186 3646 3190 3650
rect 3213 3654 3224 3657
rect 3236 3655 3244 3658
rect 3130 3639 3135 3644
rect 3139 3617 3142 3645
rect 3169 3617 3172 3641
rect 3196 3617 3199 3649
rect 3213 3648 3216 3654
rect 3236 3649 3239 3655
rect 3248 3650 3251 3653
rect 3259 3653 3262 3667
rect 3259 3650 3271 3653
rect 3259 3645 3262 3650
rect 3211 3639 3216 3644
rect 3220 3617 3223 3645
rect 3250 3617 3253 3641
rect 2867 3613 2941 3617
rect 2945 3613 2947 3617
rect 2951 3613 2955 3617
rect 2959 3613 2973 3617
rect 2977 3613 2982 3617
rect 2986 3613 2991 3617
rect 2995 3613 3014 3617
rect 3018 3613 3048 3617
rect 3052 3613 3063 3617
rect 3067 3613 3091 3617
rect 3095 3613 3108 3617
rect 3112 3613 3132 3617
rect 3136 3613 3186 3617
rect 3193 3613 3213 3617
rect 3217 3613 3267 3617
rect 2595 3597 2617 3600
rect 2621 3597 2628 3600
rect 2879 3606 2955 3610
rect 2959 3606 3014 3610
rect 3018 3606 3039 3610
rect 3043 3606 3070 3610
rect 3074 3606 3103 3610
rect 2653 3597 2677 3600
rect 2681 3597 2686 3600
rect 3002 3599 3003 3603
rect 3027 3598 3028 3602
rect 3074 3599 3075 3603
rect 2699 3594 2708 3598
rect 2586 3591 2601 3594
rect 2081 3576 2084 3580
rect 2091 3576 2094 3580
rect 2112 3576 2115 3581
rect 2139 3580 2140 3584
rect 2137 3576 2140 3580
rect 2155 3576 2158 3581
rect 2185 3580 2190 3585
rect 2194 3581 2195 3584
rect 2210 3583 2213 3589
rect 2210 3580 2218 3583
rect 2265 3580 2270 3585
rect 2274 3581 2276 3584
rect 2291 3583 2294 3589
rect 2640 3591 2659 3594
rect 2605 3587 2612 3590
rect 2637 3584 2640 3590
rect 2291 3580 2299 3583
rect 2663 3587 2670 3590
rect 2950 3585 2953 3590
rect 2957 3585 2960 3590
rect 2940 3582 2942 3585
rect 2950 3582 2960 3585
rect 2210 3577 2213 3580
rect 2291 3577 2294 3580
rect 1629 3564 1666 3568
rect 1670 3564 1696 3568
rect 1700 3564 1724 3568
rect 1728 3564 1916 3568
rect 2065 3561 2068 3565
rect 2092 3561 2093 3565
rect 2137 3561 2139 3565
rect 1629 3557 1647 3561
rect 1651 3557 1697 3561
rect 1701 3557 1748 3561
rect 1752 3557 1952 3561
rect 2010 3554 2022 3558
rect 2026 3554 2053 3558
rect 2057 3554 2075 3558
rect 2079 3554 2140 3558
rect 2144 3554 2158 3558
rect 2194 3551 2197 3569
rect 2275 3551 2278 3569
rect 2584 3568 2587 3580
rect 2605 3568 2608 3580
rect 2621 3568 2624 3580
rect 2640 3571 2652 3574
rect 2663 3568 2666 3580
rect 2679 3568 2682 3580
rect 2700 3568 2703 3580
rect 2950 3576 2953 3582
rect 2957 3576 2960 3582
rect 2966 3584 2969 3590
rect 2982 3585 2985 3590
rect 2966 3580 2968 3584
rect 2972 3580 2974 3584
rect 2982 3583 2988 3585
rect 2992 3583 2993 3585
rect 2982 3581 2993 3583
rect 3010 3583 3013 3590
rect 2966 3576 2969 3580
rect 2982 3576 2985 3581
rect 3011 3579 3013 3583
rect 3010 3576 3013 3579
rect 3026 3584 3029 3590
rect 3036 3584 3039 3590
rect 3057 3585 3060 3590
rect 3036 3580 3045 3584
rect 3057 3581 3058 3585
rect 3062 3582 3065 3585
rect 3082 3584 3085 3590
rect 3100 3585 3103 3590
rect 3139 3593 3142 3613
rect 3220 3593 3223 3613
rect 3026 3576 3029 3580
rect 3036 3576 3039 3580
rect 3057 3576 3060 3581
rect 3084 3580 3085 3584
rect 3082 3576 3085 3580
rect 3100 3576 3103 3581
rect 3130 3580 3135 3585
rect 3139 3581 3140 3584
rect 3155 3583 3158 3589
rect 3155 3580 3163 3583
rect 3210 3580 3215 3585
rect 3219 3581 3221 3584
rect 3236 3583 3239 3589
rect 3236 3580 3244 3583
rect 3155 3577 3158 3580
rect 3236 3577 3239 3580
rect 2574 3564 2611 3568
rect 2615 3564 2641 3568
rect 2645 3564 2669 3568
rect 2673 3564 2861 3568
rect 3010 3561 3013 3565
rect 3037 3561 3038 3565
rect 3082 3561 3084 3565
rect 2574 3557 2592 3561
rect 2596 3557 2642 3561
rect 2646 3557 2693 3561
rect 2697 3557 2897 3561
rect 2955 3554 2967 3558
rect 2971 3554 2998 3558
rect 3002 3554 3020 3558
rect 3024 3554 3085 3558
rect 3089 3554 3103 3558
rect 3139 3551 3142 3569
rect 3220 3551 3223 3569
rect 1910 3547 1995 3551
rect 1999 3547 2011 3551
rect 2015 3547 2029 3551
rect 2033 3547 2040 3551
rect 2044 3547 2046 3551
rect 2050 3547 2065 3551
rect 2069 3547 2102 3551
rect 2106 3547 2107 3551
rect 2111 3547 2119 3551
rect 2123 3547 2147 3551
rect 2151 3547 2163 3551
rect 2167 3547 2187 3551
rect 2191 3547 2241 3551
rect 2245 3547 2268 3551
rect 2272 3547 2330 3551
rect 2334 3547 2345 3551
rect 2855 3547 2940 3551
rect 2944 3547 2956 3551
rect 2960 3547 2974 3551
rect 2978 3547 2985 3551
rect 2989 3547 2991 3551
rect 2995 3547 3010 3551
rect 3014 3547 3047 3551
rect 3051 3547 3052 3551
rect 3056 3547 3064 3551
rect 3068 3547 3092 3551
rect 3096 3547 3108 3551
rect 3112 3547 3132 3551
rect 3136 3547 3186 3551
rect 3190 3547 3213 3551
rect 3217 3547 3275 3551
rect 3279 3547 3290 3551
rect 1946 3540 2006 3544
rect 2010 3540 2022 3544
rect 2026 3540 2053 3544
rect 2057 3540 2075 3544
rect 2079 3540 2140 3544
rect 2144 3540 2158 3544
rect 2194 3537 2197 3547
rect 2224 3543 2227 3547
rect 2275 3543 2278 3547
rect 2065 3533 2068 3537
rect 2092 3533 2093 3537
rect 2137 3533 2139 3537
rect 1994 3513 1997 3516
rect 2005 3516 2008 3522
rect 2012 3516 2015 3522
rect 2005 3513 2015 3516
rect 2005 3508 2008 3513
rect 2012 3508 2015 3513
rect 2021 3518 2024 3522
rect 2021 3514 2023 3518
rect 2027 3514 2029 3518
rect 2037 3517 2040 3522
rect 2065 3519 2068 3522
rect 2037 3515 2048 3517
rect 2021 3508 2024 3514
rect 2037 3513 2043 3515
rect 2037 3508 2040 3513
rect 2047 3513 2048 3515
rect 2066 3515 2068 3519
rect 2065 3508 2068 3515
rect 2210 3526 2213 3529
rect 2081 3518 2084 3522
rect 2091 3518 2094 3522
rect 2091 3514 2100 3518
rect 2112 3517 2115 3522
rect 2137 3518 2140 3522
rect 2081 3508 2084 3514
rect 2091 3508 2094 3514
rect 2112 3513 2113 3517
rect 2117 3513 2120 3516
rect 2139 3514 2140 3518
rect 2155 3517 2158 3522
rect 2187 3522 2198 3525
rect 2210 3523 2218 3526
rect 2112 3508 2115 3513
rect 2137 3508 2140 3514
rect 2187 3516 2190 3522
rect 2210 3517 2213 3523
rect 2222 3518 2225 3521
rect 2233 3521 2236 3535
rect 2284 3530 2287 3535
rect 2299 3537 2302 3547
rect 2329 3543 2332 3547
rect 2268 3526 2269 3529
rect 2273 3526 2276 3529
rect 2891 3540 2951 3544
rect 2955 3540 2967 3544
rect 2971 3540 2998 3544
rect 3002 3540 3020 3544
rect 3024 3540 3085 3544
rect 3089 3540 3103 3544
rect 3139 3537 3142 3547
rect 3169 3543 3172 3547
rect 3220 3543 3223 3547
rect 2315 3526 2318 3529
rect 2241 3521 2246 3526
rect 2284 3521 2287 3526
rect 2233 3518 2241 3521
rect 2155 3508 2158 3513
rect 2233 3513 2236 3518
rect 2292 3522 2303 3525
rect 2315 3523 2323 3526
rect 2185 3507 2190 3512
rect 2057 3495 2058 3499
rect 2082 3496 2083 3500
rect 2129 3495 2130 3499
rect 1934 3488 2010 3492
rect 2014 3488 2069 3492
rect 2073 3488 2094 3492
rect 2098 3488 2125 3492
rect 2129 3488 2158 3492
rect 2194 3485 2197 3513
rect 2224 3485 2227 3509
rect 2275 3485 2278 3517
rect 2292 3516 2295 3522
rect 2315 3517 2318 3523
rect 2327 3518 2330 3521
rect 2338 3521 2341 3535
rect 3010 3533 3013 3537
rect 3037 3533 3038 3537
rect 3082 3533 3084 3537
rect 2338 3518 2344 3521
rect 2338 3513 2341 3518
rect 2939 3513 2942 3516
rect 2950 3516 2953 3522
rect 2957 3516 2960 3522
rect 2950 3513 2960 3516
rect 2290 3507 2295 3512
rect 2299 3485 2302 3513
rect 2329 3485 2332 3509
rect 2950 3508 2953 3513
rect 2957 3508 2960 3513
rect 2966 3518 2969 3522
rect 2966 3514 2968 3518
rect 2972 3514 2974 3518
rect 2982 3517 2985 3522
rect 3010 3519 3013 3522
rect 2982 3515 2993 3517
rect 2966 3508 2969 3514
rect 2982 3513 2988 3515
rect 2982 3508 2985 3513
rect 2992 3513 2993 3515
rect 3011 3515 3013 3519
rect 3010 3508 3013 3515
rect 3155 3526 3158 3529
rect 3026 3518 3029 3522
rect 3036 3518 3039 3522
rect 3036 3514 3045 3518
rect 3057 3517 3060 3522
rect 3082 3518 3085 3522
rect 3026 3508 3029 3514
rect 3036 3508 3039 3514
rect 3057 3513 3058 3517
rect 3062 3513 3065 3516
rect 3084 3514 3085 3518
rect 3100 3517 3103 3522
rect 3132 3522 3143 3525
rect 3155 3523 3163 3526
rect 3057 3508 3060 3513
rect 3082 3508 3085 3514
rect 3132 3516 3135 3522
rect 3155 3517 3158 3523
rect 3167 3518 3170 3521
rect 3178 3521 3181 3535
rect 3229 3530 3232 3535
rect 3244 3537 3247 3547
rect 3274 3543 3277 3547
rect 3213 3526 3214 3529
rect 3218 3526 3221 3529
rect 3260 3526 3263 3529
rect 3186 3521 3191 3526
rect 3229 3521 3232 3526
rect 3178 3518 3186 3521
rect 3100 3508 3103 3513
rect 3178 3513 3181 3518
rect 3237 3522 3248 3525
rect 3260 3523 3268 3526
rect 3130 3507 3135 3512
rect 3002 3495 3003 3499
rect 3027 3496 3028 3500
rect 3074 3495 3075 3499
rect 2879 3488 2955 3492
rect 2959 3488 3014 3492
rect 3018 3488 3039 3492
rect 3043 3488 3070 3492
rect 3074 3488 3103 3492
rect 3139 3485 3142 3513
rect 3169 3485 3172 3509
rect 3220 3485 3223 3517
rect 3237 3516 3240 3522
rect 3260 3517 3263 3523
rect 3272 3518 3275 3521
rect 3283 3521 3286 3535
rect 3283 3518 3289 3521
rect 3283 3513 3286 3518
rect 3235 3507 3240 3512
rect 3244 3485 3247 3513
rect 3274 3485 3277 3509
rect 1922 3481 1996 3485
rect 2000 3481 2002 3485
rect 2006 3481 2010 3485
rect 2014 3481 2028 3485
rect 2032 3481 2037 3485
rect 2041 3481 2046 3485
rect 2050 3481 2069 3485
rect 2073 3481 2103 3485
rect 2107 3481 2118 3485
rect 2122 3481 2146 3485
rect 2150 3481 2163 3485
rect 2167 3481 2187 3485
rect 2191 3481 2241 3485
rect 2245 3481 2268 3485
rect 2272 3481 2292 3485
rect 2296 3481 2344 3485
rect 2867 3481 2941 3485
rect 2945 3481 2947 3485
rect 2951 3481 2955 3485
rect 2959 3481 2973 3485
rect 2977 3481 2982 3485
rect 2986 3481 2991 3485
rect 2995 3481 3014 3485
rect 3018 3481 3048 3485
rect 3052 3481 3063 3485
rect 3067 3481 3091 3485
rect 3095 3481 3108 3485
rect 3112 3481 3132 3485
rect 3136 3481 3186 3485
rect 3190 3481 3213 3485
rect 3217 3481 3237 3485
rect 3241 3481 3289 3485
rect 1934 3474 2010 3478
rect 2014 3474 2069 3478
rect 2073 3474 2094 3478
rect 2098 3474 2125 3478
rect 2129 3474 2158 3478
rect 2057 3467 2058 3471
rect 2082 3466 2083 3470
rect 2129 3467 2130 3471
rect 2194 3462 2197 3481
rect 2299 3462 2302 3481
rect 2879 3474 2955 3478
rect 2959 3474 3014 3478
rect 3018 3474 3039 3478
rect 3043 3474 3070 3478
rect 3074 3474 3103 3478
rect 3002 3467 3003 3471
rect 3027 3466 3028 3470
rect 3074 3467 3075 3471
rect 3139 3462 3142 3481
rect 3244 3462 3247 3481
rect 2005 3453 2008 3458
rect 2012 3453 2015 3458
rect 1995 3450 1997 3453
rect 2005 3450 2015 3453
rect 2005 3444 2008 3450
rect 2012 3444 2015 3450
rect 2021 3452 2024 3458
rect 2037 3453 2040 3458
rect 2021 3448 2023 3452
rect 2027 3448 2029 3452
rect 2037 3451 2043 3453
rect 2047 3451 2048 3453
rect 2037 3449 2048 3451
rect 2065 3451 2068 3458
rect 2021 3444 2024 3448
rect 2037 3444 2040 3449
rect 2066 3447 2068 3451
rect 2065 3444 2068 3447
rect 2081 3452 2084 3458
rect 2091 3452 2094 3458
rect 2112 3453 2115 3458
rect 2091 3448 2100 3452
rect 2112 3449 2113 3453
rect 2117 3450 2120 3453
rect 2137 3452 2140 3458
rect 2155 3453 2158 3458
rect 2081 3444 2084 3448
rect 2091 3444 2094 3448
rect 2112 3444 2115 3449
rect 2139 3448 2140 3452
rect 2184 3449 2189 3454
rect 2193 3450 2195 3453
rect 2210 3452 2213 3458
rect 2210 3449 2218 3452
rect 2290 3449 2295 3454
rect 2299 3450 2300 3453
rect 2315 3452 2318 3458
rect 2315 3449 2323 3452
rect 2950 3453 2953 3458
rect 2957 3453 2960 3458
rect 2940 3450 2942 3453
rect 2950 3450 2960 3453
rect 2137 3444 2140 3448
rect 2155 3444 2158 3449
rect 2210 3446 2213 3449
rect 2315 3446 2318 3449
rect 2950 3444 2953 3450
rect 2065 3429 2068 3433
rect 2092 3429 2093 3433
rect 2137 3429 2139 3433
rect 1946 3422 2022 3426
rect 2026 3422 2053 3426
rect 2057 3422 2075 3426
rect 2079 3422 2140 3426
rect 2144 3422 2158 3426
rect 2194 3419 2197 3438
rect 2299 3419 2302 3438
rect 2957 3444 2960 3450
rect 2966 3452 2969 3458
rect 2982 3453 2985 3458
rect 2966 3448 2968 3452
rect 2972 3448 2974 3452
rect 2982 3451 2988 3453
rect 2992 3451 2993 3453
rect 2982 3449 2993 3451
rect 3010 3451 3013 3458
rect 2966 3444 2969 3448
rect 2982 3444 2985 3449
rect 3011 3447 3013 3451
rect 3010 3444 3013 3447
rect 3026 3452 3029 3458
rect 3036 3452 3039 3458
rect 3057 3453 3060 3458
rect 3036 3448 3045 3452
rect 3057 3449 3058 3453
rect 3062 3450 3065 3453
rect 3082 3452 3085 3458
rect 3100 3453 3103 3458
rect 3026 3444 3029 3448
rect 3036 3444 3039 3448
rect 3057 3444 3060 3449
rect 3084 3448 3085 3452
rect 3129 3449 3134 3454
rect 3138 3450 3140 3453
rect 3155 3452 3158 3458
rect 3155 3449 3163 3452
rect 3235 3449 3240 3454
rect 3244 3450 3245 3453
rect 3260 3452 3263 3458
rect 3260 3449 3268 3452
rect 3082 3444 3085 3448
rect 3100 3444 3103 3449
rect 3155 3446 3158 3449
rect 3260 3446 3263 3449
rect 3010 3429 3013 3433
rect 3037 3429 3038 3433
rect 3082 3429 3084 3433
rect 2891 3422 2967 3426
rect 2971 3422 2998 3426
rect 3002 3422 3020 3426
rect 3024 3422 3085 3426
rect 3089 3422 3103 3426
rect 3139 3419 3142 3438
rect 3244 3419 3247 3438
rect 1910 3415 1995 3419
rect 1999 3415 2011 3419
rect 2015 3415 2029 3419
rect 2033 3415 2040 3419
rect 2044 3415 2046 3419
rect 2050 3415 2065 3419
rect 2069 3415 2102 3419
rect 2106 3415 2107 3419
rect 2111 3415 2119 3419
rect 2123 3415 2147 3419
rect 2151 3415 2163 3419
rect 2167 3415 2187 3419
rect 2191 3415 2241 3419
rect 2245 3415 2268 3419
rect 2272 3415 2322 3419
rect 2326 3415 2330 3419
rect 2334 3415 2358 3419
rect 2362 3415 2412 3419
rect 2855 3415 2940 3419
rect 2944 3415 2956 3419
rect 2960 3415 2974 3419
rect 2978 3415 2985 3419
rect 2989 3415 2991 3419
rect 2995 3415 3010 3419
rect 3014 3415 3047 3419
rect 3051 3415 3052 3419
rect 3056 3415 3064 3419
rect 3068 3415 3092 3419
rect 3096 3415 3108 3419
rect 3112 3415 3132 3419
rect 3136 3415 3186 3419
rect 3190 3415 3213 3419
rect 3217 3415 3267 3419
rect 3271 3415 3275 3419
rect 3279 3415 3303 3419
rect 3307 3415 3357 3419
rect 1946 3408 2022 3412
rect 2026 3408 2053 3412
rect 2057 3408 2075 3412
rect 2079 3408 2140 3412
rect 2144 3408 2158 3412
rect 2194 3405 2197 3415
rect 2224 3411 2227 3415
rect 2251 3411 2254 3415
rect 2065 3401 2068 3405
rect 2092 3401 2093 3405
rect 2137 3401 2139 3405
rect 1994 3381 1997 3384
rect 2005 3384 2008 3390
rect 2012 3384 2015 3390
rect 2005 3381 2015 3384
rect 2005 3376 2008 3381
rect 2012 3376 2015 3381
rect 2021 3386 2024 3390
rect 2021 3382 2023 3386
rect 2027 3382 2029 3386
rect 2037 3385 2040 3390
rect 2065 3387 2068 3390
rect 2037 3383 2048 3385
rect 2021 3376 2024 3382
rect 2037 3381 2043 3383
rect 2037 3376 2040 3381
rect 2047 3381 2048 3383
rect 2066 3383 2068 3387
rect 2065 3376 2068 3383
rect 2210 3394 2213 3397
rect 2081 3386 2084 3390
rect 2091 3386 2094 3390
rect 2091 3382 2100 3386
rect 2112 3385 2115 3390
rect 2137 3386 2140 3390
rect 2081 3376 2084 3382
rect 2091 3376 2094 3382
rect 2112 3381 2113 3385
rect 2117 3381 2120 3384
rect 2139 3382 2140 3386
rect 2155 3385 2158 3390
rect 2187 3390 2198 3393
rect 2210 3391 2218 3394
rect 2112 3376 2115 3381
rect 2137 3376 2140 3382
rect 2187 3384 2190 3390
rect 2210 3385 2213 3391
rect 2222 3386 2225 3389
rect 2233 3389 2236 3403
rect 2260 3398 2263 3403
rect 2275 3405 2278 3415
rect 2305 3411 2308 3415
rect 2341 3411 2344 3415
rect 2244 3394 2245 3397
rect 2249 3394 2252 3397
rect 2291 3394 2294 3397
rect 2233 3386 2241 3389
rect 2260 3389 2263 3394
rect 2155 3376 2158 3381
rect 2233 3381 2236 3386
rect 2241 3382 2245 3386
rect 2268 3390 2279 3393
rect 2291 3391 2299 3394
rect 2185 3375 2190 3380
rect 2057 3363 2058 3367
rect 2082 3364 2083 3368
rect 2129 3363 2130 3367
rect 1934 3356 2010 3360
rect 2014 3356 2069 3360
rect 2073 3356 2094 3360
rect 2098 3356 2125 3360
rect 2129 3356 2158 3360
rect 2194 3353 2197 3381
rect 2224 3353 2227 3377
rect 2251 3353 2254 3385
rect 2268 3384 2271 3390
rect 2291 3385 2294 3391
rect 2303 3386 2306 3389
rect 2314 3389 2317 3403
rect 2350 3398 2353 3403
rect 2365 3405 2368 3415
rect 2395 3411 2398 3415
rect 2339 3394 2342 3397
rect 2891 3408 2967 3412
rect 2971 3408 2998 3412
rect 3002 3408 3020 3412
rect 3024 3408 3085 3412
rect 3089 3408 3103 3412
rect 3139 3405 3142 3415
rect 3169 3411 3172 3415
rect 3196 3411 3199 3415
rect 2381 3394 2384 3397
rect 2314 3386 2323 3389
rect 2350 3389 2353 3394
rect 2314 3381 2317 3386
rect 2266 3375 2271 3380
rect 2275 3353 2278 3381
rect 2357 3392 2369 3393
rect 2361 3390 2369 3392
rect 2381 3391 2389 3394
rect 2381 3385 2384 3391
rect 2393 3386 2396 3389
rect 2404 3389 2407 3403
rect 3010 3401 3013 3405
rect 3037 3401 3038 3405
rect 3082 3401 3084 3405
rect 2404 3386 2424 3389
rect 2305 3353 2308 3377
rect 2341 3353 2344 3385
rect 2404 3381 2407 3386
rect 2939 3381 2942 3384
rect 2950 3384 2953 3390
rect 2957 3384 2960 3390
rect 2950 3381 2960 3384
rect 2365 3353 2368 3381
rect 2395 3353 2398 3377
rect 2950 3376 2953 3381
rect 2957 3376 2960 3381
rect 2966 3386 2969 3390
rect 2966 3382 2968 3386
rect 2972 3382 2974 3386
rect 2982 3385 2985 3390
rect 3010 3387 3013 3390
rect 2982 3383 2993 3385
rect 2966 3376 2969 3382
rect 2982 3381 2988 3383
rect 2982 3376 2985 3381
rect 2992 3381 2993 3383
rect 3011 3383 3013 3387
rect 3010 3376 3013 3383
rect 3155 3394 3158 3397
rect 3026 3386 3029 3390
rect 3036 3386 3039 3390
rect 3036 3382 3045 3386
rect 3057 3385 3060 3390
rect 3082 3386 3085 3390
rect 3026 3376 3029 3382
rect 3036 3376 3039 3382
rect 3057 3381 3058 3385
rect 3062 3381 3065 3384
rect 3084 3382 3085 3386
rect 3100 3385 3103 3390
rect 3132 3390 3143 3393
rect 3155 3391 3163 3394
rect 3057 3376 3060 3381
rect 3082 3376 3085 3382
rect 3132 3384 3135 3390
rect 3155 3385 3158 3391
rect 3167 3386 3170 3389
rect 3178 3389 3181 3403
rect 3205 3398 3208 3403
rect 3220 3405 3223 3415
rect 3250 3411 3253 3415
rect 3286 3411 3289 3415
rect 3189 3394 3190 3397
rect 3194 3394 3197 3397
rect 3236 3394 3239 3397
rect 3178 3386 3186 3389
rect 3205 3389 3208 3394
rect 3100 3376 3103 3381
rect 3178 3381 3181 3386
rect 3186 3382 3190 3386
rect 3213 3390 3224 3393
rect 3236 3391 3244 3394
rect 3130 3375 3135 3380
rect 3002 3363 3003 3367
rect 3027 3364 3028 3368
rect 3074 3363 3075 3367
rect 2879 3356 2955 3360
rect 2959 3356 3014 3360
rect 3018 3356 3039 3360
rect 3043 3356 3070 3360
rect 3074 3356 3103 3360
rect 3139 3353 3142 3381
rect 3169 3353 3172 3377
rect 3196 3353 3199 3385
rect 3213 3384 3216 3390
rect 3236 3385 3239 3391
rect 3248 3386 3251 3389
rect 3259 3389 3262 3403
rect 3295 3398 3298 3403
rect 3310 3405 3313 3415
rect 3340 3411 3343 3415
rect 3284 3394 3287 3397
rect 3326 3394 3329 3397
rect 3259 3386 3268 3389
rect 3295 3389 3298 3394
rect 3259 3381 3262 3386
rect 3211 3375 3216 3380
rect 3220 3353 3223 3381
rect 3302 3392 3314 3393
rect 3306 3390 3314 3392
rect 3326 3391 3334 3394
rect 3326 3385 3329 3391
rect 3338 3386 3341 3389
rect 3349 3389 3352 3403
rect 3349 3386 3369 3389
rect 3250 3353 3253 3377
rect 3286 3353 3289 3385
rect 3349 3381 3352 3386
rect 3310 3353 3313 3381
rect 3340 3353 3343 3377
rect 1922 3349 1996 3353
rect 2000 3349 2002 3353
rect 2006 3349 2010 3353
rect 2014 3349 2028 3353
rect 2032 3349 2037 3353
rect 2041 3349 2046 3353
rect 2050 3349 2069 3353
rect 2073 3349 2103 3353
rect 2107 3349 2118 3353
rect 2122 3349 2146 3353
rect 2150 3349 2163 3353
rect 2167 3349 2187 3353
rect 2191 3349 2241 3353
rect 2248 3349 2268 3353
rect 2272 3349 2322 3353
rect 2326 3349 2358 3353
rect 2362 3349 2412 3353
rect 2867 3349 2941 3353
rect 2945 3349 2947 3353
rect 2951 3349 2955 3353
rect 2959 3349 2973 3353
rect 2977 3349 2982 3353
rect 2986 3349 2991 3353
rect 2995 3349 3014 3353
rect 3018 3349 3048 3353
rect 3052 3349 3063 3353
rect 3067 3349 3091 3353
rect 3095 3349 3108 3353
rect 3112 3349 3132 3353
rect 3136 3349 3186 3353
rect 3193 3349 3213 3353
rect 3217 3349 3267 3353
rect 3271 3349 3303 3353
rect 3307 3349 3357 3353
rect 1934 3342 2010 3346
rect 2014 3342 2069 3346
rect 2073 3342 2094 3346
rect 2098 3342 2125 3346
rect 2129 3342 2158 3346
rect 2057 3335 2058 3339
rect 2082 3334 2083 3338
rect 2129 3335 2130 3339
rect 2005 3321 2008 3326
rect 2012 3321 2015 3326
rect 1995 3318 1997 3321
rect 2005 3318 2015 3321
rect 2005 3312 2008 3318
rect 2012 3312 2015 3318
rect 2021 3320 2024 3326
rect 2037 3321 2040 3326
rect 2021 3316 2023 3320
rect 2027 3316 2029 3320
rect 2037 3319 2043 3321
rect 2047 3319 2048 3321
rect 2037 3317 2048 3319
rect 2065 3319 2068 3326
rect 2021 3312 2024 3316
rect 2037 3312 2040 3317
rect 2066 3315 2068 3319
rect 2065 3312 2068 3315
rect 2081 3320 2084 3326
rect 2091 3320 2094 3326
rect 2112 3321 2115 3326
rect 2091 3316 2100 3320
rect 2112 3317 2113 3321
rect 2117 3318 2120 3321
rect 2137 3320 2140 3326
rect 2155 3321 2158 3326
rect 2194 3327 2197 3349
rect 2275 3327 2278 3349
rect 2365 3327 2368 3349
rect 2879 3342 2955 3346
rect 2959 3342 3014 3346
rect 3018 3342 3039 3346
rect 3043 3342 3070 3346
rect 3074 3342 3103 3346
rect 3002 3335 3003 3339
rect 3027 3334 3028 3338
rect 3074 3335 3075 3339
rect 2081 3312 2084 3316
rect 2091 3312 2094 3316
rect 2112 3312 2115 3317
rect 2139 3316 2140 3320
rect 2137 3312 2140 3316
rect 2155 3312 2158 3317
rect 2185 3314 2190 3319
rect 2194 3315 2195 3318
rect 2210 3317 2213 3323
rect 2210 3314 2218 3317
rect 2265 3314 2270 3319
rect 2274 3315 2276 3318
rect 2291 3317 2294 3323
rect 2291 3314 2299 3317
rect 2358 3315 2366 3318
rect 2381 3317 2384 3323
rect 2950 3321 2953 3326
rect 2957 3321 2960 3326
rect 2940 3318 2942 3321
rect 2381 3314 2389 3317
rect 2950 3318 2960 3321
rect 2210 3311 2213 3314
rect 2291 3311 2294 3314
rect 2381 3311 2384 3314
rect 2950 3312 2953 3318
rect 2065 3297 2068 3301
rect 2092 3297 2093 3301
rect 2137 3297 2139 3301
rect 2957 3312 2960 3318
rect 2966 3320 2969 3326
rect 2982 3321 2985 3326
rect 2966 3316 2968 3320
rect 2972 3316 2974 3320
rect 2982 3319 2988 3321
rect 2992 3319 2993 3321
rect 2982 3317 2993 3319
rect 3010 3319 3013 3326
rect 2966 3312 2969 3316
rect 2982 3312 2985 3317
rect 3011 3315 3013 3319
rect 3010 3312 3013 3315
rect 3026 3320 3029 3326
rect 3036 3320 3039 3326
rect 3057 3321 3060 3326
rect 3036 3316 3045 3320
rect 3057 3317 3058 3321
rect 3062 3318 3065 3321
rect 3082 3320 3085 3326
rect 3100 3321 3103 3326
rect 3139 3327 3142 3349
rect 3220 3327 3223 3349
rect 3310 3327 3313 3349
rect 3026 3312 3029 3316
rect 3036 3312 3039 3316
rect 3057 3312 3060 3317
rect 3084 3316 3085 3320
rect 3082 3312 3085 3316
rect 3100 3312 3103 3317
rect 3130 3314 3135 3319
rect 3139 3315 3140 3318
rect 3155 3317 3158 3323
rect 3155 3314 3163 3317
rect 3210 3314 3215 3319
rect 3219 3315 3221 3318
rect 3236 3317 3239 3323
rect 3236 3314 3244 3317
rect 3303 3315 3311 3318
rect 3326 3317 3329 3323
rect 3326 3314 3334 3317
rect 3155 3311 3158 3314
rect 3236 3311 3239 3314
rect 3326 3311 3329 3314
rect 1946 3290 2022 3294
rect 2026 3290 2053 3294
rect 2057 3290 2075 3294
rect 2079 3290 2140 3294
rect 2144 3290 2158 3294
rect 2194 3287 2197 3303
rect 2275 3287 2278 3303
rect 2365 3287 2368 3303
rect 3010 3297 3013 3301
rect 3037 3297 3038 3301
rect 3082 3297 3084 3301
rect 2891 3290 2967 3294
rect 2971 3290 2998 3294
rect 3002 3290 3020 3294
rect 3024 3290 3085 3294
rect 3089 3290 3103 3294
rect 3139 3287 3142 3303
rect 3220 3287 3223 3303
rect 3310 3287 3313 3303
rect 1910 3283 1995 3287
rect 1999 3283 2011 3287
rect 2015 3283 2029 3287
rect 2033 3283 2040 3287
rect 2044 3283 2046 3287
rect 2050 3283 2065 3287
rect 2069 3283 2102 3287
rect 2106 3283 2107 3287
rect 2111 3283 2119 3287
rect 2123 3283 2147 3287
rect 2151 3283 2163 3287
rect 2167 3283 2187 3287
rect 2191 3283 2241 3287
rect 2245 3283 2268 3287
rect 2272 3283 2358 3287
rect 2362 3283 2416 3287
rect 2855 3283 2940 3287
rect 2944 3283 2956 3287
rect 2960 3283 2974 3287
rect 2978 3283 2985 3287
rect 2989 3283 2991 3287
rect 2995 3283 3010 3287
rect 3014 3283 3047 3287
rect 3051 3283 3052 3287
rect 3056 3283 3064 3287
rect 3068 3283 3092 3287
rect 3096 3283 3108 3287
rect 3112 3283 3132 3287
rect 3136 3283 3186 3287
rect 3190 3283 3213 3287
rect 3217 3283 3303 3287
rect 3307 3283 3361 3287
rect 1946 3276 2022 3280
rect 2026 3276 2053 3280
rect 2057 3276 2075 3280
rect 2079 3276 2140 3280
rect 2144 3276 2158 3280
rect 2194 3273 2197 3283
rect 2224 3279 2227 3283
rect 2065 3269 2068 3273
rect 2092 3269 2093 3273
rect 2137 3269 2139 3273
rect 1994 3249 1997 3252
rect 2005 3252 2008 3258
rect 2012 3252 2015 3258
rect 2005 3249 2015 3252
rect 2005 3244 2008 3249
rect 2012 3244 2015 3249
rect 2021 3254 2024 3258
rect 2021 3250 2023 3254
rect 2027 3250 2029 3254
rect 2037 3253 2040 3258
rect 2065 3255 2068 3258
rect 2037 3251 2048 3253
rect 2021 3244 2024 3250
rect 2037 3249 2043 3251
rect 2037 3244 2040 3249
rect 2047 3249 2048 3251
rect 2066 3251 2068 3255
rect 2065 3244 2068 3251
rect 2891 3276 2967 3280
rect 2971 3276 2998 3280
rect 3002 3276 3020 3280
rect 3024 3276 3085 3280
rect 3089 3276 3103 3280
rect 3139 3273 3142 3283
rect 3169 3279 3172 3283
rect 2210 3262 2213 3265
rect 2081 3254 2084 3258
rect 2091 3254 2094 3258
rect 2091 3250 2100 3254
rect 2112 3253 2115 3258
rect 2137 3254 2140 3258
rect 2081 3244 2084 3250
rect 2091 3244 2094 3250
rect 2112 3249 2113 3253
rect 2117 3249 2120 3252
rect 2139 3250 2140 3254
rect 2155 3253 2158 3258
rect 2187 3258 2198 3261
rect 2210 3259 2218 3262
rect 2112 3244 2115 3249
rect 2137 3244 2140 3250
rect 2187 3252 2190 3258
rect 2210 3253 2213 3259
rect 2222 3254 2225 3257
rect 2233 3257 2236 3271
rect 3010 3269 3013 3273
rect 3037 3269 3038 3273
rect 3082 3269 3084 3273
rect 2241 3257 2246 3262
rect 2233 3254 2241 3257
rect 2155 3244 2158 3249
rect 2233 3249 2236 3254
rect 2939 3249 2942 3252
rect 2950 3252 2953 3258
rect 2957 3252 2960 3258
rect 2950 3249 2960 3252
rect 2185 3243 2190 3248
rect 1495 3235 1616 3239
rect 1504 3228 1513 3232
rect 1517 3228 1549 3232
rect 1553 3228 1616 3232
rect 1620 3228 1645 3232
rect 1649 3228 1681 3232
rect 1685 3228 1748 3232
rect 1752 3228 1777 3232
rect 1781 3228 1813 3232
rect 1817 3228 1880 3232
rect 1884 3228 1964 3232
rect 2057 3231 2058 3235
rect 2082 3232 2083 3236
rect 2129 3231 2130 3235
rect 1504 3221 1537 3225
rect 1541 3221 1565 3225
rect 1569 3221 1595 3225
rect 1599 3221 1632 3225
rect 1636 3221 1669 3225
rect 1673 3221 1697 3225
rect 1701 3221 1727 3225
rect 1731 3221 1764 3225
rect 1768 3221 1801 3225
rect 1805 3221 1829 3225
rect 1833 3221 1859 3225
rect 1863 3221 1896 3225
rect 1900 3221 1904 3225
rect 1989 3224 2010 3228
rect 2014 3224 2019 3228
rect 2023 3224 2069 3228
rect 2073 3224 2094 3228
rect 2098 3224 2125 3228
rect 2129 3224 2158 3228
rect 2194 3221 2197 3249
rect 2224 3221 2227 3245
rect 2950 3244 2953 3249
rect 2957 3244 2960 3249
rect 2966 3254 2969 3258
rect 2966 3250 2968 3254
rect 2972 3250 2974 3254
rect 2982 3253 2985 3258
rect 3010 3255 3013 3258
rect 2982 3251 2993 3253
rect 2966 3244 2969 3250
rect 2982 3249 2988 3251
rect 2982 3244 2985 3249
rect 2992 3249 2993 3251
rect 3011 3251 3013 3255
rect 3010 3244 3013 3251
rect 3155 3262 3158 3265
rect 3026 3254 3029 3258
rect 3036 3254 3039 3258
rect 3036 3250 3045 3254
rect 3057 3253 3060 3258
rect 3082 3254 3085 3258
rect 3026 3244 3029 3250
rect 3036 3244 3039 3250
rect 3057 3249 3058 3253
rect 3062 3249 3065 3252
rect 3084 3250 3085 3254
rect 3100 3253 3103 3258
rect 3132 3258 3143 3261
rect 3155 3259 3163 3262
rect 3057 3244 3060 3249
rect 3082 3244 3085 3250
rect 3132 3252 3135 3258
rect 3155 3253 3158 3259
rect 3167 3254 3170 3257
rect 3178 3257 3181 3271
rect 3186 3257 3191 3262
rect 3178 3254 3186 3257
rect 3100 3244 3103 3249
rect 3178 3249 3181 3254
rect 3130 3243 3135 3248
rect 2449 3228 2458 3232
rect 2462 3228 2494 3232
rect 2498 3228 2561 3232
rect 2565 3228 2590 3232
rect 2594 3228 2626 3232
rect 2630 3228 2693 3232
rect 2697 3228 2722 3232
rect 2726 3228 2758 3232
rect 2762 3228 2825 3232
rect 2829 3228 2909 3232
rect 3002 3231 3003 3235
rect 3027 3232 3028 3236
rect 3074 3231 3075 3235
rect 2449 3221 2482 3225
rect 2486 3221 2510 3225
rect 2514 3221 2540 3225
rect 2544 3221 2577 3225
rect 2581 3221 2614 3225
rect 2618 3221 2642 3225
rect 2646 3221 2672 3225
rect 2676 3221 2709 3225
rect 2713 3221 2746 3225
rect 2750 3221 2774 3225
rect 2778 3221 2804 3225
rect 2808 3221 2841 3225
rect 2845 3221 2849 3225
rect 2934 3224 2955 3228
rect 2959 3224 2964 3228
rect 2968 3224 3014 3228
rect 3018 3224 3039 3228
rect 3043 3224 3070 3228
rect 3074 3224 3103 3228
rect 3139 3221 3142 3249
rect 3169 3221 3172 3245
rect 1507 3211 1510 3221
rect 1528 3211 1531 3221
rect 1544 3211 1547 3221
rect 1558 3214 1563 3218
rect 1567 3214 1574 3218
rect 1586 3211 1589 3221
rect 1602 3211 1605 3221
rect 1623 3211 1626 3221
rect 1639 3211 1642 3221
rect 1660 3211 1663 3221
rect 1676 3211 1679 3221
rect 1690 3214 1695 3218
rect 1699 3214 1706 3218
rect 1718 3211 1721 3221
rect 1734 3211 1737 3221
rect 1755 3211 1758 3221
rect 1771 3211 1774 3221
rect 1792 3211 1795 3221
rect 1808 3211 1811 3221
rect 1822 3214 1827 3218
rect 1831 3214 1838 3218
rect 1850 3211 1853 3221
rect 1866 3211 1869 3221
rect 1887 3211 1890 3221
rect 1922 3217 1996 3221
rect 2000 3217 2002 3221
rect 2006 3217 2010 3221
rect 2014 3217 2028 3221
rect 2032 3217 2037 3221
rect 2041 3217 2046 3221
rect 2050 3217 2069 3221
rect 2073 3217 2103 3221
rect 2107 3217 2118 3221
rect 2122 3217 2146 3221
rect 2150 3217 2163 3221
rect 2167 3217 2187 3221
rect 2191 3217 2271 3221
rect 2275 3217 2289 3221
rect 2293 3217 2298 3221
rect 2302 3217 2307 3221
rect 2311 3217 2330 3221
rect 2334 3217 2364 3221
rect 2368 3217 2379 3221
rect 2383 3217 2407 3221
rect 2411 3217 2420 3221
rect 1524 3197 1529 3200
rect 1533 3197 1557 3200
rect 1582 3197 1589 3200
rect 1593 3197 1615 3200
rect 1635 3197 1642 3200
rect 1656 3197 1661 3200
rect 1665 3197 1689 3200
rect 1714 3197 1721 3200
rect 1725 3197 1747 3200
rect 1767 3197 1774 3200
rect 1788 3197 1793 3200
rect 1797 3197 1821 3200
rect 1934 3210 2010 3214
rect 2014 3210 2019 3214
rect 2023 3210 2069 3214
rect 2073 3210 2094 3214
rect 2098 3210 2125 3214
rect 2129 3210 2158 3214
rect 1846 3197 1853 3200
rect 1857 3197 1879 3200
rect 2057 3203 2058 3207
rect 2082 3202 2083 3206
rect 2129 3203 2130 3207
rect 1540 3187 1547 3190
rect 1551 3191 1570 3194
rect 1570 3184 1573 3190
rect 1598 3187 1605 3190
rect 1609 3191 1624 3194
rect 1672 3187 1679 3190
rect 1683 3191 1702 3194
rect 1702 3184 1705 3190
rect 1730 3187 1737 3190
rect 1741 3191 1756 3194
rect 1804 3187 1811 3190
rect 1815 3191 1834 3194
rect 1834 3184 1837 3190
rect 1862 3187 1869 3190
rect 1873 3191 1890 3194
rect 2005 3189 2008 3194
rect 2012 3189 2015 3194
rect 1995 3186 1997 3189
rect 2005 3186 2015 3189
rect 2005 3180 2008 3186
rect 1507 3168 1510 3180
rect 1528 3168 1531 3180
rect 1544 3168 1547 3180
rect 1558 3171 1570 3174
rect 1586 3168 1589 3180
rect 1602 3168 1605 3180
rect 1623 3168 1626 3180
rect 1639 3168 1642 3180
rect 1660 3168 1663 3180
rect 1676 3168 1679 3180
rect 1690 3171 1702 3174
rect 1718 3168 1721 3180
rect 1734 3168 1737 3180
rect 1755 3168 1758 3180
rect 1771 3168 1774 3180
rect 1792 3168 1795 3180
rect 1808 3168 1811 3180
rect 1822 3171 1834 3174
rect 1850 3168 1853 3180
rect 1866 3168 1869 3180
rect 1887 3168 1890 3180
rect 2012 3180 2015 3186
rect 2021 3188 2024 3194
rect 2037 3189 2040 3194
rect 2021 3184 2023 3188
rect 2027 3184 2029 3188
rect 2037 3187 2043 3189
rect 2047 3187 2048 3189
rect 2037 3185 2048 3187
rect 2065 3187 2068 3194
rect 2021 3180 2024 3184
rect 2037 3180 2040 3185
rect 2066 3183 2068 3187
rect 2065 3180 2068 3183
rect 2081 3188 2084 3194
rect 2091 3188 2094 3194
rect 2112 3189 2115 3194
rect 2091 3184 2100 3188
rect 2112 3185 2113 3189
rect 2117 3186 2120 3189
rect 2137 3188 2140 3194
rect 2155 3189 2158 3194
rect 2194 3191 2197 3217
rect 2230 3210 2249 3214
rect 2253 3210 2271 3214
rect 2275 3210 2330 3214
rect 2334 3210 2355 3214
rect 2359 3210 2386 3214
rect 2390 3210 2419 3214
rect 2452 3211 2455 3221
rect 2473 3211 2476 3221
rect 2489 3211 2492 3221
rect 2503 3214 2508 3218
rect 2512 3214 2519 3218
rect 2531 3211 2534 3221
rect 2547 3211 2550 3221
rect 2568 3211 2571 3221
rect 2584 3211 2587 3221
rect 2605 3211 2608 3221
rect 2621 3211 2624 3221
rect 2635 3214 2640 3218
rect 2644 3214 2651 3218
rect 2663 3211 2666 3221
rect 2679 3211 2682 3221
rect 2700 3211 2703 3221
rect 2716 3211 2719 3221
rect 2737 3211 2740 3221
rect 2753 3211 2756 3221
rect 2767 3214 2772 3218
rect 2776 3214 2783 3218
rect 2795 3211 2798 3221
rect 2811 3211 2814 3221
rect 2832 3211 2835 3221
rect 2867 3217 2941 3221
rect 2945 3217 2947 3221
rect 2951 3217 2955 3221
rect 2959 3217 2973 3221
rect 2977 3217 2982 3221
rect 2986 3217 2991 3221
rect 2995 3217 3014 3221
rect 3018 3217 3048 3221
rect 3052 3217 3063 3221
rect 3067 3217 3091 3221
rect 3095 3217 3108 3221
rect 3112 3217 3132 3221
rect 3136 3217 3216 3221
rect 3220 3217 3234 3221
rect 3238 3217 3243 3221
rect 3247 3217 3252 3221
rect 3256 3217 3275 3221
rect 3279 3217 3309 3221
rect 3313 3217 3324 3221
rect 3328 3217 3352 3221
rect 3356 3217 3365 3221
rect 2230 3198 2233 3210
rect 2318 3203 2319 3207
rect 2343 3202 2344 3206
rect 2390 3203 2391 3207
rect 2081 3180 2084 3184
rect 2091 3180 2094 3184
rect 2112 3180 2115 3185
rect 2139 3184 2140 3188
rect 2257 3189 2260 3194
rect 2266 3189 2269 3194
rect 2273 3189 2276 3194
rect 2137 3180 2140 3184
rect 2155 3180 2158 3185
rect 2184 3178 2189 3183
rect 2193 3179 2195 3182
rect 2210 3181 2213 3187
rect 2242 3186 2276 3189
rect 2210 3178 2218 3181
rect 2210 3175 2213 3178
rect 1504 3164 1537 3168
rect 1541 3164 1565 3168
rect 1569 3164 1595 3168
rect 1599 3164 1669 3168
rect 1673 3164 1697 3168
rect 1701 3164 1727 3168
rect 1731 3164 1801 3168
rect 1805 3164 1829 3168
rect 1833 3164 1859 3168
rect 1863 3164 1916 3168
rect 2065 3165 2068 3169
rect 2092 3165 2093 3169
rect 2137 3165 2139 3169
rect 2242 3172 2245 3186
rect 2266 3180 2269 3186
rect 2273 3180 2276 3186
rect 2282 3188 2285 3194
rect 2298 3189 2301 3194
rect 2282 3184 2284 3188
rect 2288 3184 2290 3188
rect 2298 3187 2304 3189
rect 2308 3187 2309 3189
rect 2298 3185 2309 3187
rect 2326 3187 2329 3194
rect 2282 3180 2285 3184
rect 2298 3180 2301 3185
rect 2327 3183 2329 3187
rect 2326 3180 2329 3183
rect 2469 3197 2474 3200
rect 2478 3197 2502 3200
rect 2527 3197 2534 3200
rect 2538 3197 2560 3200
rect 2580 3197 2587 3200
rect 2601 3197 2606 3200
rect 2610 3197 2634 3200
rect 2659 3197 2666 3200
rect 2670 3197 2692 3200
rect 2712 3197 2719 3200
rect 2733 3197 2738 3200
rect 2742 3197 2766 3200
rect 2879 3210 2955 3214
rect 2959 3210 2964 3214
rect 2968 3210 3014 3214
rect 3018 3210 3039 3214
rect 3043 3210 3070 3214
rect 3074 3210 3103 3214
rect 2791 3197 2798 3200
rect 2802 3197 2824 3200
rect 3002 3203 3003 3207
rect 3027 3202 3028 3206
rect 3074 3203 3075 3207
rect 2342 3188 2345 3194
rect 2352 3188 2355 3194
rect 2373 3189 2376 3194
rect 2352 3184 2361 3188
rect 2373 3185 2374 3189
rect 2378 3186 2381 3189
rect 2398 3188 2401 3194
rect 2416 3189 2419 3194
rect 2342 3180 2345 3184
rect 2352 3180 2355 3184
rect 2373 3180 2376 3185
rect 2400 3184 2401 3188
rect 2398 3180 2401 3184
rect 2416 3180 2419 3185
rect 2485 3187 2492 3190
rect 2496 3191 2515 3194
rect 2515 3184 2518 3190
rect 2543 3187 2550 3190
rect 2554 3191 2569 3194
rect 2617 3187 2624 3190
rect 2628 3191 2647 3194
rect 2647 3184 2650 3190
rect 2675 3187 2682 3190
rect 2686 3191 2701 3194
rect 2749 3187 2756 3190
rect 2760 3191 2779 3194
rect 2779 3184 2782 3190
rect 2807 3187 2814 3190
rect 2818 3191 2835 3194
rect 2950 3189 2953 3194
rect 2957 3189 2960 3194
rect 2940 3186 2942 3189
rect 2950 3186 2960 3189
rect 2950 3180 2953 3186
rect 1504 3157 1513 3161
rect 1517 3157 1564 3161
rect 1568 3157 1614 3161
rect 1618 3157 1645 3161
rect 1649 3157 1696 3161
rect 1700 3157 1746 3161
rect 1750 3157 1777 3161
rect 1781 3157 1828 3161
rect 1832 3157 1878 3161
rect 1882 3158 1952 3161
rect 2008 3158 2022 3162
rect 2026 3158 2053 3162
rect 2057 3158 2075 3162
rect 2079 3158 2140 3162
rect 2144 3158 2158 3162
rect 2194 3155 2197 3167
rect 2326 3165 2329 3169
rect 2353 3165 2354 3169
rect 2398 3165 2400 3169
rect 2452 3168 2455 3180
rect 2473 3168 2476 3180
rect 2489 3168 2492 3180
rect 2503 3171 2515 3174
rect 2531 3168 2534 3180
rect 2547 3168 2550 3180
rect 2568 3168 2571 3180
rect 2584 3168 2587 3180
rect 2605 3168 2608 3180
rect 2621 3168 2624 3180
rect 2635 3171 2647 3174
rect 2663 3168 2666 3180
rect 2679 3168 2682 3180
rect 2700 3168 2703 3180
rect 2716 3168 2719 3180
rect 2737 3168 2740 3180
rect 2753 3168 2756 3180
rect 2767 3171 2779 3174
rect 2795 3168 2798 3180
rect 2811 3168 2814 3180
rect 2832 3168 2835 3180
rect 2957 3180 2960 3186
rect 2966 3188 2969 3194
rect 2982 3189 2985 3194
rect 2966 3184 2968 3188
rect 2972 3184 2974 3188
rect 2982 3187 2988 3189
rect 2992 3187 2993 3189
rect 2982 3185 2993 3187
rect 3010 3187 3013 3194
rect 2966 3180 2969 3184
rect 2982 3180 2985 3185
rect 3011 3183 3013 3187
rect 3010 3180 3013 3183
rect 3026 3188 3029 3194
rect 3036 3188 3039 3194
rect 3057 3189 3060 3194
rect 3036 3184 3045 3188
rect 3057 3185 3058 3189
rect 3062 3186 3065 3189
rect 3082 3188 3085 3194
rect 3100 3189 3103 3194
rect 3139 3191 3142 3217
rect 3175 3210 3194 3214
rect 3198 3210 3216 3214
rect 3220 3210 3275 3214
rect 3279 3210 3300 3214
rect 3304 3210 3331 3214
rect 3335 3210 3364 3214
rect 3175 3198 3178 3210
rect 3263 3203 3264 3207
rect 3288 3202 3289 3206
rect 3335 3203 3336 3207
rect 3026 3180 3029 3184
rect 3036 3180 3039 3184
rect 3057 3180 3060 3185
rect 3084 3184 3085 3188
rect 3202 3189 3205 3194
rect 3211 3189 3214 3194
rect 3218 3189 3221 3194
rect 3082 3180 3085 3184
rect 3100 3180 3103 3185
rect 3129 3178 3134 3183
rect 3138 3179 3140 3182
rect 3155 3181 3158 3187
rect 3187 3186 3221 3189
rect 3155 3178 3163 3181
rect 3155 3175 3158 3178
rect 2449 3164 2482 3168
rect 2486 3164 2510 3168
rect 2514 3164 2540 3168
rect 2544 3164 2614 3168
rect 2618 3164 2642 3168
rect 2646 3164 2672 3168
rect 2676 3164 2746 3168
rect 2750 3164 2774 3168
rect 2778 3164 2804 3168
rect 2808 3164 2861 3168
rect 3010 3165 3013 3169
rect 3037 3165 3038 3169
rect 3082 3165 3084 3169
rect 3187 3172 3190 3186
rect 3211 3180 3214 3186
rect 3218 3180 3221 3186
rect 3227 3188 3230 3194
rect 3243 3189 3246 3194
rect 3227 3184 3229 3188
rect 3233 3184 3235 3188
rect 3243 3187 3249 3189
rect 3253 3187 3254 3189
rect 3243 3185 3254 3187
rect 3271 3187 3274 3194
rect 3227 3180 3230 3184
rect 3243 3180 3246 3185
rect 3272 3183 3274 3187
rect 3271 3180 3274 3183
rect 3287 3188 3290 3194
rect 3297 3188 3300 3194
rect 3318 3189 3321 3194
rect 3297 3184 3306 3188
rect 3318 3185 3319 3189
rect 3323 3186 3326 3189
rect 3343 3188 3346 3194
rect 3361 3189 3364 3194
rect 3287 3180 3290 3184
rect 3297 3180 3300 3184
rect 3318 3180 3321 3185
rect 3345 3184 3346 3188
rect 3343 3180 3346 3184
rect 3361 3180 3364 3185
rect 2234 3158 2239 3162
rect 2243 3158 2283 3162
rect 2287 3158 2314 3162
rect 2318 3158 2336 3162
rect 2340 3158 2401 3162
rect 2405 3158 2419 3162
rect 2449 3157 2458 3161
rect 2462 3157 2509 3161
rect 2513 3157 2559 3161
rect 2563 3157 2590 3161
rect 2594 3157 2641 3161
rect 2645 3157 2691 3161
rect 2695 3157 2722 3161
rect 2726 3157 2773 3161
rect 2777 3157 2823 3161
rect 2827 3158 2897 3161
rect 2953 3158 2967 3162
rect 2971 3158 2998 3162
rect 3002 3158 3020 3162
rect 3024 3158 3085 3162
rect 3089 3158 3103 3162
rect 3139 3155 3142 3167
rect 3271 3165 3274 3169
rect 3298 3165 3299 3169
rect 3343 3165 3345 3169
rect 3179 3158 3184 3162
rect 3188 3158 3228 3162
rect 3232 3158 3259 3162
rect 3263 3158 3281 3162
rect 3285 3158 3346 3162
rect 3350 3158 3364 3162
rect 1511 3151 1895 3154
rect 1910 3151 1995 3155
rect 1999 3151 2011 3155
rect 2015 3151 2029 3155
rect 2033 3151 2040 3155
rect 2044 3151 2046 3155
rect 2050 3151 2065 3155
rect 2069 3151 2102 3155
rect 2106 3151 2107 3155
rect 2111 3151 2119 3155
rect 2123 3151 2147 3155
rect 2151 3151 2187 3155
rect 2191 3151 2230 3155
rect 2234 3151 2241 3155
rect 2245 3151 2256 3155
rect 2260 3151 2272 3155
rect 2276 3151 2290 3155
rect 2294 3151 2301 3155
rect 2305 3151 2307 3155
rect 2311 3151 2326 3155
rect 2330 3151 2363 3155
rect 2367 3151 2368 3155
rect 2372 3151 2380 3155
rect 2384 3151 2408 3155
rect 2412 3151 2420 3155
rect 2456 3151 2840 3154
rect 2855 3151 2940 3155
rect 2944 3151 2956 3155
rect 2960 3151 2974 3155
rect 2978 3151 2985 3155
rect 2989 3151 2991 3155
rect 2995 3151 3010 3155
rect 3014 3151 3047 3155
rect 3051 3151 3052 3155
rect 3056 3151 3064 3155
rect 3068 3151 3092 3155
rect 3096 3151 3132 3155
rect 3136 3151 3175 3155
rect 3179 3151 3186 3155
rect 3190 3151 3201 3155
rect 3205 3151 3217 3155
rect 3221 3151 3235 3155
rect 3239 3151 3246 3155
rect 3250 3151 3252 3155
rect 3256 3151 3271 3155
rect 3275 3151 3308 3155
rect 3312 3151 3313 3155
rect 3317 3151 3325 3155
rect 3329 3151 3353 3155
rect 3357 3151 3365 3155
rect 1654 3144 1763 3147
rect 1946 3144 2004 3148
rect 2008 3144 2238 3147
rect 2428 3145 2436 3149
rect 2599 3144 2708 3147
rect 2891 3144 2949 3148
rect 2953 3144 3183 3147
rect 3373 3145 3381 3149
rect 1634 3136 1638 3140
rect 1642 3136 1646 3140
rect 1934 3137 2248 3140
rect 1622 3135 1626 3136
rect 1654 3135 1658 3136
rect 1982 3130 2255 3133
rect 2424 3127 2428 3132
rect 2579 3136 2583 3140
rect 2587 3136 2591 3140
rect 2879 3137 3193 3140
rect 2567 3135 2571 3136
rect 2599 3135 2603 3136
rect 2927 3130 3198 3134
rect 3369 3127 3373 3132
rect 1495 3123 1622 3127
rect 1626 3123 1642 3127
rect 1658 3123 2567 3127
rect 2571 3123 2587 3127
rect 2603 3123 3461 3127
rect 1650 3116 1895 3119
rect 1970 3116 2296 3120
rect 2300 3116 2332 3120
rect 2336 3116 2399 3120
rect 2403 3116 2419 3120
rect 2595 3116 2840 3119
rect 2915 3116 3241 3120
rect 3245 3116 3277 3120
rect 3281 3116 3344 3120
rect 3348 3116 3364 3120
rect 1665 3109 1895 3112
rect 1910 3109 2282 3113
rect 2286 3109 2320 3113
rect 2324 3109 2348 3113
rect 2352 3109 2378 3113
rect 2382 3109 2415 3113
rect 1634 3100 1638 3104
rect 1642 3100 1646 3104
rect 2290 3099 2293 3109
rect 2311 3099 2314 3109
rect 2327 3099 2330 3109
rect 2341 3102 2346 3106
rect 2350 3102 2357 3106
rect 2369 3099 2372 3109
rect 2385 3099 2388 3109
rect 2406 3099 2409 3109
rect 2610 3109 2840 3112
rect 2855 3109 3227 3113
rect 3231 3109 3265 3113
rect 3269 3109 3293 3113
rect 3297 3109 3323 3113
rect 3327 3109 3360 3113
rect 2579 3100 2583 3104
rect 2587 3100 2591 3104
rect 3235 3099 3238 3109
rect 3256 3099 3259 3109
rect 3272 3099 3275 3109
rect 3286 3102 3291 3106
rect 3295 3102 3302 3106
rect 3314 3099 3317 3109
rect 3330 3099 3333 3109
rect 3351 3099 3354 3109
rect 1654 3093 1764 3096
rect 1504 3086 1513 3090
rect 1517 3086 1549 3090
rect 1553 3086 1616 3090
rect 1620 3086 1645 3090
rect 1649 3086 1681 3090
rect 1685 3086 1748 3090
rect 1752 3086 1777 3090
rect 1781 3086 1813 3090
rect 1817 3086 1880 3090
rect 1884 3086 1964 3090
rect 1504 3079 1537 3083
rect 1541 3079 1565 3083
rect 1569 3079 1595 3083
rect 1599 3079 1632 3083
rect 1636 3079 1669 3083
rect 1673 3079 1697 3083
rect 1701 3079 1727 3083
rect 1731 3079 1764 3083
rect 1768 3079 1801 3083
rect 1805 3079 1829 3083
rect 1833 3079 1859 3083
rect 1863 3079 1896 3083
rect 1900 3079 1904 3083
rect 2307 3085 2312 3088
rect 2316 3085 2340 3088
rect 2599 3093 2709 3096
rect 2365 3085 2372 3088
rect 2376 3085 2398 3088
rect 2449 3086 2458 3090
rect 2462 3086 2494 3090
rect 2498 3086 2561 3090
rect 2565 3086 2590 3090
rect 2594 3086 2626 3090
rect 2630 3086 2693 3090
rect 2697 3086 2722 3090
rect 2726 3086 2758 3090
rect 2762 3086 2825 3090
rect 2829 3086 2909 3090
rect 1507 3069 1510 3079
rect 1528 3069 1531 3079
rect 1544 3069 1547 3079
rect 1558 3072 1563 3076
rect 1567 3072 1574 3076
rect 1586 3069 1589 3079
rect 1602 3069 1605 3079
rect 1623 3069 1626 3079
rect 1639 3069 1642 3079
rect 1660 3069 1663 3079
rect 1676 3069 1679 3079
rect 1690 3072 1695 3076
rect 1699 3072 1706 3076
rect 1718 3069 1721 3079
rect 1734 3069 1737 3079
rect 1755 3069 1758 3079
rect 1771 3069 1774 3079
rect 1792 3069 1795 3079
rect 1808 3069 1811 3079
rect 1822 3072 1827 3076
rect 1831 3072 1838 3076
rect 1850 3069 1853 3079
rect 1866 3069 1869 3079
rect 1887 3069 1890 3079
rect 2323 3075 2330 3078
rect 2334 3079 2353 3082
rect 1524 3055 1529 3058
rect 1533 3055 1557 3058
rect 1582 3055 1589 3058
rect 1593 3055 1615 3058
rect 1635 3055 1642 3058
rect 1656 3055 1661 3058
rect 1665 3055 1689 3058
rect 1714 3055 1721 3058
rect 1725 3055 1747 3058
rect 1767 3055 1774 3058
rect 1788 3055 1793 3058
rect 1797 3055 1821 3058
rect 1846 3055 1853 3058
rect 1857 3055 1879 3058
rect 2353 3072 2356 3078
rect 2381 3075 2388 3078
rect 2392 3079 2407 3082
rect 2449 3079 2482 3083
rect 2486 3079 2510 3083
rect 2514 3079 2540 3083
rect 2544 3079 2577 3083
rect 2581 3079 2614 3083
rect 2618 3079 2642 3083
rect 2646 3079 2672 3083
rect 2676 3079 2709 3083
rect 2713 3079 2746 3083
rect 2750 3079 2774 3083
rect 2778 3079 2804 3083
rect 2808 3079 2841 3083
rect 2845 3079 2849 3083
rect 3252 3085 3257 3088
rect 3261 3085 3285 3088
rect 3310 3085 3317 3088
rect 3321 3085 3343 3088
rect 2452 3069 2455 3079
rect 2473 3069 2476 3079
rect 2489 3069 2492 3079
rect 2503 3072 2508 3076
rect 2512 3072 2519 3076
rect 2531 3069 2534 3079
rect 2547 3069 2550 3079
rect 2568 3069 2571 3079
rect 2584 3069 2587 3079
rect 2605 3069 2608 3079
rect 2621 3069 2624 3079
rect 2635 3072 2640 3076
rect 2644 3072 2651 3076
rect 2663 3069 2666 3079
rect 2679 3069 2682 3079
rect 2700 3069 2703 3079
rect 2716 3069 2719 3079
rect 2737 3069 2740 3079
rect 2753 3069 2756 3079
rect 2767 3072 2772 3076
rect 2776 3072 2783 3076
rect 2795 3069 2798 3079
rect 2811 3069 2814 3079
rect 2832 3069 2835 3079
rect 3268 3075 3275 3078
rect 3279 3079 3298 3082
rect 2290 3056 2293 3068
rect 2311 3056 2314 3068
rect 2327 3056 2330 3068
rect 2341 3059 2353 3062
rect 2369 3056 2372 3068
rect 2385 3056 2388 3068
rect 2406 3056 2409 3068
rect 1540 3045 1547 3048
rect 1551 3049 1570 3052
rect 1570 3042 1573 3048
rect 1598 3045 1605 3048
rect 1609 3049 1624 3052
rect 1672 3045 1679 3048
rect 1683 3049 1702 3052
rect 1702 3042 1705 3048
rect 1730 3045 1737 3048
rect 1741 3049 1756 3052
rect 1804 3045 1811 3048
rect 1815 3049 1834 3052
rect 1834 3042 1837 3048
rect 1862 3045 1869 3048
rect 1873 3049 1890 3052
rect 1922 3052 2320 3056
rect 2324 3052 2348 3056
rect 2352 3052 2378 3056
rect 2382 3052 2419 3056
rect 2469 3055 2474 3058
rect 2478 3055 2502 3058
rect 2527 3055 2534 3058
rect 2538 3055 2560 3058
rect 2580 3055 2587 3058
rect 2601 3055 2606 3058
rect 2610 3055 2634 3058
rect 2659 3055 2666 3058
rect 2670 3055 2692 3058
rect 2712 3055 2719 3058
rect 2733 3055 2738 3058
rect 2742 3055 2766 3058
rect 2791 3055 2798 3058
rect 2802 3055 2824 3058
rect 3298 3072 3301 3078
rect 3326 3075 3333 3078
rect 3337 3079 3352 3082
rect 3235 3056 3238 3068
rect 3256 3056 3259 3068
rect 3272 3056 3275 3068
rect 3286 3059 3298 3062
rect 3314 3056 3317 3068
rect 3330 3056 3333 3068
rect 3351 3056 3354 3068
rect 1958 3045 2296 3049
rect 2300 3045 2347 3049
rect 2351 3045 2397 3049
rect 2401 3045 2419 3049
rect 2485 3045 2492 3048
rect 2496 3049 2515 3052
rect 1507 3026 1510 3038
rect 1528 3026 1531 3038
rect 1544 3026 1547 3038
rect 1558 3029 1570 3032
rect 1586 3026 1589 3038
rect 1602 3026 1605 3038
rect 1623 3026 1626 3038
rect 1639 3026 1642 3038
rect 1660 3026 1663 3038
rect 1676 3026 1679 3038
rect 1690 3029 1702 3032
rect 1718 3026 1721 3038
rect 1734 3026 1737 3038
rect 1755 3026 1758 3038
rect 1771 3026 1774 3038
rect 1792 3026 1795 3038
rect 1808 3026 1811 3038
rect 1822 3029 1834 3032
rect 1850 3026 1853 3038
rect 1866 3026 1869 3038
rect 1887 3026 1890 3038
rect 2293 3038 2414 3041
rect 2515 3042 2518 3048
rect 2543 3045 2550 3048
rect 2554 3049 2569 3052
rect 2617 3045 2624 3048
rect 2628 3049 2647 3052
rect 2647 3042 2650 3048
rect 2675 3045 2682 3048
rect 2686 3049 2701 3052
rect 2749 3045 2756 3048
rect 2760 3049 2779 3052
rect 2779 3042 2782 3048
rect 2807 3045 2814 3048
rect 2818 3049 2835 3052
rect 2867 3052 3265 3056
rect 3269 3052 3293 3056
rect 3297 3052 3323 3056
rect 3327 3052 3364 3056
rect 2903 3045 3241 3049
rect 3245 3045 3292 3049
rect 3296 3045 3342 3049
rect 3346 3045 3364 3049
rect 1970 3030 2296 3034
rect 2300 3030 2332 3034
rect 2336 3030 2399 3034
rect 2403 3030 2419 3034
rect 1504 3022 1537 3026
rect 1541 3022 1565 3026
rect 1569 3022 1595 3026
rect 1599 3022 1669 3026
rect 1673 3022 1697 3026
rect 1701 3022 1727 3026
rect 1731 3022 1801 3026
rect 1805 3022 1829 3026
rect 1833 3022 1859 3026
rect 1863 3022 1916 3026
rect 2286 3023 2320 3027
rect 2324 3023 2348 3027
rect 2352 3023 2378 3027
rect 2382 3023 2415 3027
rect 2452 3026 2455 3038
rect 2473 3026 2476 3038
rect 2489 3026 2492 3038
rect 2503 3029 2515 3032
rect 2531 3026 2534 3038
rect 2547 3026 2550 3038
rect 2568 3026 2571 3038
rect 2584 3026 2587 3038
rect 2605 3026 2608 3038
rect 2621 3026 2624 3038
rect 2635 3029 2647 3032
rect 2663 3026 2666 3038
rect 2679 3026 2682 3038
rect 2700 3026 2703 3038
rect 2716 3026 2719 3038
rect 2737 3026 2740 3038
rect 2753 3026 2756 3038
rect 2767 3029 2779 3032
rect 2795 3026 2798 3038
rect 2811 3026 2814 3038
rect 2832 3026 2835 3038
rect 3238 3038 3359 3041
rect 2915 3030 3241 3034
rect 3245 3030 3277 3034
rect 3281 3030 3344 3034
rect 3348 3030 3364 3034
rect 1504 3015 1513 3019
rect 1517 3015 1564 3019
rect 1568 3015 1614 3019
rect 1618 3015 1645 3019
rect 1649 3015 1696 3019
rect 1700 3015 1746 3019
rect 1750 3015 1777 3019
rect 1781 3015 1828 3019
rect 1832 3015 1878 3019
rect 1882 3015 1952 3019
rect 2290 3013 2293 3023
rect 2311 3013 2314 3023
rect 2327 3013 2330 3023
rect 2341 3016 2346 3020
rect 2350 3016 2357 3020
rect 2369 3013 2372 3023
rect 2385 3013 2388 3023
rect 2406 3013 2409 3023
rect 2449 3022 2482 3026
rect 2486 3022 2510 3026
rect 2514 3022 2540 3026
rect 2544 3022 2614 3026
rect 2618 3022 2642 3026
rect 2646 3022 2672 3026
rect 2676 3022 2746 3026
rect 2750 3022 2774 3026
rect 2778 3022 2804 3026
rect 2808 3022 2861 3026
rect 3231 3023 3265 3027
rect 3269 3023 3293 3027
rect 3297 3023 3323 3027
rect 3327 3023 3360 3027
rect 2449 3015 2458 3019
rect 2462 3015 2509 3019
rect 2513 3015 2559 3019
rect 2563 3015 2590 3019
rect 2594 3015 2641 3019
rect 2645 3015 2691 3019
rect 2695 3015 2722 3019
rect 2726 3015 2773 3019
rect 2777 3015 2823 3019
rect 2827 3015 2897 3019
rect 3235 3013 3238 3023
rect 3256 3013 3259 3023
rect 3272 3013 3275 3023
rect 3286 3016 3291 3020
rect 3295 3016 3302 3020
rect 3314 3013 3317 3023
rect 3330 3013 3333 3023
rect 3351 3013 3354 3023
rect 1510 3008 1895 3011
rect 1504 3000 1513 3004
rect 1517 3000 1549 3004
rect 1553 3000 1616 3004
rect 1620 3000 1645 3004
rect 1649 3000 1681 3004
rect 1685 3000 1748 3004
rect 1752 3000 1777 3004
rect 1781 3000 1813 3004
rect 1817 3000 1880 3004
rect 1884 3000 1964 3004
rect 1504 2993 1537 2997
rect 1541 2993 1565 2997
rect 1569 2993 1595 2997
rect 1599 2993 1632 2997
rect 1636 2993 1669 2997
rect 1673 2993 1697 2997
rect 1701 2993 1727 2997
rect 1731 2993 1764 2997
rect 1768 2993 1801 2997
rect 1805 2993 1829 2997
rect 1833 2993 1859 2997
rect 1863 2993 1896 2997
rect 1900 2993 1904 2997
rect 2307 2999 2312 3002
rect 2316 2999 2340 3002
rect 2455 3008 2840 3011
rect 2365 2999 2372 3002
rect 2376 2999 2398 3002
rect 2449 3000 2458 3004
rect 2462 3000 2494 3004
rect 2498 3000 2561 3004
rect 2565 3000 2590 3004
rect 2594 3000 2626 3004
rect 2630 3000 2693 3004
rect 2697 3000 2722 3004
rect 2726 3000 2758 3004
rect 2762 3000 2825 3004
rect 2829 3000 2909 3004
rect 1507 2983 1510 2993
rect 1528 2983 1531 2993
rect 1544 2983 1547 2993
rect 1558 2986 1563 2990
rect 1567 2986 1574 2990
rect 1586 2983 1589 2993
rect 1602 2983 1605 2993
rect 1623 2983 1626 2993
rect 1639 2983 1642 2993
rect 1660 2983 1663 2993
rect 1676 2983 1679 2993
rect 1690 2986 1695 2990
rect 1699 2986 1706 2990
rect 1718 2983 1721 2993
rect 1734 2983 1737 2993
rect 1755 2983 1758 2993
rect 1771 2983 1774 2993
rect 1792 2983 1795 2993
rect 1808 2983 1811 2993
rect 1822 2986 1827 2990
rect 1831 2986 1838 2990
rect 1850 2983 1853 2993
rect 1866 2983 1869 2993
rect 1887 2983 1890 2993
rect 2323 2989 2330 2992
rect 2334 2993 2353 2996
rect 1524 2969 1529 2972
rect 1533 2969 1557 2972
rect 1582 2969 1589 2972
rect 1593 2969 1615 2972
rect 1635 2969 1642 2972
rect 1656 2969 1661 2972
rect 1665 2969 1689 2972
rect 1714 2969 1721 2972
rect 1725 2969 1747 2972
rect 1767 2969 1774 2972
rect 1788 2969 1793 2972
rect 1797 2969 1821 2972
rect 1846 2969 1853 2972
rect 1857 2969 1879 2972
rect 2353 2986 2356 2992
rect 2381 2989 2388 2992
rect 2392 2993 2407 2996
rect 2418 2991 2429 2995
rect 2449 2993 2482 2997
rect 2486 2993 2510 2997
rect 2514 2993 2540 2997
rect 2544 2993 2577 2997
rect 2581 2993 2614 2997
rect 2618 2993 2642 2997
rect 2646 2993 2672 2997
rect 2676 2993 2709 2997
rect 2713 2993 2746 2997
rect 2750 2993 2774 2997
rect 2778 2993 2804 2997
rect 2808 2993 2841 2997
rect 2845 2993 2849 2997
rect 3252 2999 3257 3002
rect 3261 2999 3285 3002
rect 3310 2999 3317 3002
rect 3321 2999 3343 3002
rect 2452 2983 2455 2993
rect 2473 2983 2476 2993
rect 2489 2983 2492 2993
rect 2503 2986 2508 2990
rect 2512 2986 2519 2990
rect 2531 2983 2534 2993
rect 2547 2983 2550 2993
rect 2568 2983 2571 2993
rect 2584 2983 2587 2993
rect 2605 2983 2608 2993
rect 2621 2983 2624 2993
rect 2635 2986 2640 2990
rect 2644 2986 2651 2990
rect 2663 2983 2666 2993
rect 2679 2983 2682 2993
rect 2700 2983 2703 2993
rect 2716 2983 2719 2993
rect 2737 2983 2740 2993
rect 2753 2983 2756 2993
rect 2767 2986 2772 2990
rect 2776 2986 2783 2990
rect 2795 2983 2798 2993
rect 2811 2983 2814 2993
rect 2832 2983 2835 2993
rect 3268 2989 3275 2992
rect 3279 2993 3298 2996
rect 2290 2970 2293 2982
rect 2311 2970 2314 2982
rect 2327 2970 2330 2982
rect 2341 2973 2353 2976
rect 2369 2970 2372 2982
rect 2385 2970 2388 2982
rect 2406 2970 2409 2982
rect 1540 2959 1547 2962
rect 1551 2963 1570 2966
rect 1570 2956 1573 2962
rect 1598 2959 1605 2962
rect 1609 2963 1624 2966
rect 1672 2959 1679 2962
rect 1683 2963 1702 2966
rect 1702 2956 1705 2962
rect 1730 2959 1737 2962
rect 1741 2963 1756 2966
rect 1804 2959 1811 2962
rect 1815 2963 1834 2966
rect 1834 2956 1837 2962
rect 1862 2959 1869 2962
rect 1873 2963 1890 2966
rect 1922 2966 2320 2970
rect 2324 2966 2348 2970
rect 2352 2966 2378 2970
rect 2382 2966 2419 2970
rect 2469 2969 2474 2972
rect 2478 2969 2502 2972
rect 2527 2969 2534 2972
rect 2538 2969 2560 2972
rect 2580 2969 2587 2972
rect 2601 2969 2606 2972
rect 2610 2969 2634 2972
rect 2659 2969 2666 2972
rect 2670 2969 2692 2972
rect 2712 2969 2719 2972
rect 2733 2969 2738 2972
rect 2742 2969 2766 2972
rect 2791 2969 2798 2972
rect 2802 2969 2824 2972
rect 3298 2986 3301 2992
rect 3326 2989 3333 2992
rect 3337 2993 3352 2996
rect 3363 2991 3374 2995
rect 3235 2970 3238 2982
rect 3256 2970 3259 2982
rect 3272 2970 3275 2982
rect 3286 2973 3298 2976
rect 3314 2970 3317 2982
rect 3330 2970 3333 2982
rect 3351 2970 3354 2982
rect 1958 2959 2296 2963
rect 2300 2959 2347 2963
rect 2351 2959 2397 2963
rect 2401 2959 2419 2963
rect 2485 2959 2492 2962
rect 2496 2963 2515 2966
rect 2515 2956 2518 2962
rect 2543 2959 2550 2962
rect 2554 2963 2569 2966
rect 2617 2959 2624 2962
rect 2628 2963 2647 2966
rect 2647 2956 2650 2962
rect 2675 2959 2682 2962
rect 2686 2963 2701 2966
rect 2749 2959 2756 2962
rect 2760 2963 2779 2966
rect 2779 2956 2782 2962
rect 2807 2959 2814 2962
rect 2818 2963 2835 2966
rect 2867 2966 3265 2970
rect 3269 2966 3293 2970
rect 3297 2966 3323 2970
rect 3327 2966 3364 2970
rect 2903 2959 3241 2963
rect 3245 2959 3292 2963
rect 3296 2959 3342 2963
rect 3346 2959 3364 2963
rect 1507 2940 1510 2952
rect 1528 2940 1531 2952
rect 1544 2940 1547 2952
rect 1558 2943 1570 2946
rect 1586 2940 1589 2952
rect 1602 2940 1605 2952
rect 1623 2940 1626 2952
rect 1639 2940 1642 2952
rect 1660 2940 1663 2952
rect 1676 2940 1679 2952
rect 1690 2943 1702 2946
rect 1718 2940 1721 2952
rect 1734 2940 1737 2952
rect 1755 2940 1758 2952
rect 1771 2940 1774 2952
rect 1792 2940 1795 2952
rect 1808 2940 1811 2952
rect 1822 2943 1834 2946
rect 1850 2940 1853 2952
rect 1866 2940 1869 2952
rect 1887 2940 1890 2952
rect 2452 2940 2455 2952
rect 2473 2940 2476 2952
rect 2489 2940 2492 2952
rect 2503 2943 2515 2946
rect 2531 2940 2534 2952
rect 2547 2940 2550 2952
rect 2568 2940 2571 2952
rect 2584 2940 2587 2952
rect 2605 2940 2608 2952
rect 2621 2940 2624 2952
rect 2635 2943 2647 2946
rect 2663 2940 2666 2952
rect 2679 2940 2682 2952
rect 2700 2940 2703 2952
rect 2716 2940 2719 2952
rect 2737 2940 2740 2952
rect 2753 2940 2756 2952
rect 2767 2943 2779 2946
rect 2795 2940 2798 2952
rect 2811 2940 2814 2952
rect 2832 2940 2835 2952
rect 1504 2936 1537 2940
rect 1541 2936 1565 2940
rect 1569 2936 1595 2940
rect 1599 2936 1669 2940
rect 1673 2936 1697 2940
rect 1701 2936 1727 2940
rect 1731 2936 1801 2940
rect 1805 2936 1829 2940
rect 1833 2936 1859 2940
rect 1863 2936 1916 2940
rect 2449 2936 2482 2940
rect 2486 2936 2510 2940
rect 2514 2936 2540 2940
rect 2544 2936 2614 2940
rect 2618 2936 2642 2940
rect 2646 2936 2672 2940
rect 2676 2936 2746 2940
rect 2750 2936 2774 2940
rect 2778 2936 2804 2940
rect 2808 2936 2861 2940
rect 1504 2929 1513 2933
rect 1517 2929 1564 2933
rect 1568 2929 1614 2933
rect 1618 2929 1645 2933
rect 1649 2929 1696 2933
rect 1700 2929 1746 2933
rect 1750 2929 1777 2933
rect 1781 2929 1828 2933
rect 1832 2929 1878 2933
rect 1882 2929 1952 2933
rect 2449 2929 2458 2933
rect 2462 2929 2509 2933
rect 2513 2929 2559 2933
rect 2563 2929 2590 2933
rect 2594 2929 2641 2933
rect 2645 2929 2691 2933
rect 2695 2929 2722 2933
rect 2726 2929 2773 2933
rect 2777 2929 2823 2933
rect 2827 2929 2897 2933
rect 1510 2923 1895 2926
rect 2455 2923 2840 2926
rect 1635 2916 1739 2919
rect 2580 2916 2684 2919
rect 1751 2908 1755 2912
rect 1759 2908 1763 2912
rect 2696 2908 2700 2912
rect 2704 2908 2708 2912
rect 1494 2897 1739 2901
rect 1743 2897 1759 2901
rect 1775 2897 2436 2901
rect 2440 2897 2684 2901
rect 2688 2897 2704 2901
rect 2720 2897 3381 2901
rect 3385 2897 3463 2901
rect 1767 2890 1895 2893
rect 2712 2890 2840 2893
rect 1782 2883 1895 2886
rect 2727 2883 2840 2886
rect 1751 2874 1755 2878
rect 1759 2874 1763 2878
rect 2696 2874 2700 2878
rect 2704 2874 2708 2878
rect 1635 2867 1739 2870
rect 2580 2867 2684 2870
rect 1504 2860 1513 2864
rect 1517 2860 1549 2864
rect 1553 2860 1616 2864
rect 1620 2860 1645 2864
rect 1649 2860 1681 2864
rect 1685 2860 1748 2864
rect 1752 2860 1777 2864
rect 1781 2860 1813 2864
rect 1817 2860 1880 2864
rect 1884 2860 1964 2864
rect 2449 2860 2458 2864
rect 2462 2860 2494 2864
rect 2498 2860 2561 2864
rect 2565 2860 2590 2864
rect 2594 2860 2626 2864
rect 2630 2860 2693 2864
rect 2697 2860 2722 2864
rect 2726 2860 2758 2864
rect 2762 2860 2825 2864
rect 2829 2860 2909 2864
rect 1504 2853 1537 2857
rect 1541 2853 1565 2857
rect 1569 2853 1595 2857
rect 1599 2853 1632 2857
rect 1636 2853 1669 2857
rect 1673 2853 1697 2857
rect 1701 2853 1727 2857
rect 1731 2853 1764 2857
rect 1768 2853 1801 2857
rect 1805 2853 1829 2857
rect 1833 2853 1859 2857
rect 1863 2853 1896 2857
rect 1900 2853 1904 2857
rect 2449 2853 2482 2857
rect 2486 2853 2510 2857
rect 2514 2853 2540 2857
rect 2544 2853 2577 2857
rect 2581 2853 2614 2857
rect 2618 2853 2642 2857
rect 2646 2853 2672 2857
rect 2676 2853 2709 2857
rect 2713 2853 2746 2857
rect 2750 2853 2774 2857
rect 2778 2853 2804 2857
rect 2808 2853 2841 2857
rect 2845 2853 2849 2857
rect 1507 2843 1510 2853
rect 1528 2843 1531 2853
rect 1544 2843 1547 2853
rect 1558 2846 1563 2850
rect 1567 2846 1574 2850
rect 1586 2843 1589 2853
rect 1602 2843 1605 2853
rect 1623 2843 1626 2853
rect 1639 2843 1642 2853
rect 1660 2843 1663 2853
rect 1676 2843 1679 2853
rect 1690 2846 1695 2850
rect 1699 2846 1706 2850
rect 1718 2843 1721 2853
rect 1734 2843 1737 2853
rect 1755 2843 1758 2853
rect 1771 2843 1774 2853
rect 1792 2843 1795 2853
rect 1808 2843 1811 2853
rect 1822 2846 1827 2850
rect 1831 2846 1838 2850
rect 1850 2843 1853 2853
rect 1866 2843 1869 2853
rect 1887 2843 1890 2853
rect 2452 2843 2455 2853
rect 2473 2843 2476 2853
rect 2489 2843 2492 2853
rect 2503 2846 2508 2850
rect 2512 2846 2519 2850
rect 2531 2843 2534 2853
rect 2547 2843 2550 2853
rect 2568 2843 2571 2853
rect 2584 2843 2587 2853
rect 2605 2843 2608 2853
rect 2621 2843 2624 2853
rect 2635 2846 2640 2850
rect 2644 2846 2651 2850
rect 2663 2843 2666 2853
rect 2679 2843 2682 2853
rect 2700 2843 2703 2853
rect 2716 2843 2719 2853
rect 2737 2843 2740 2853
rect 2753 2843 2756 2853
rect 2767 2846 2772 2850
rect 2776 2846 2783 2850
rect 2795 2843 2798 2853
rect 2811 2843 2814 2853
rect 2832 2843 2835 2853
rect 1524 2829 1529 2832
rect 1533 2829 1557 2832
rect 1582 2829 1589 2832
rect 1593 2829 1615 2832
rect 1635 2829 1642 2832
rect 1656 2829 1661 2832
rect 1665 2829 1689 2832
rect 1714 2829 1721 2832
rect 1725 2829 1747 2832
rect 1767 2829 1774 2832
rect 1788 2829 1793 2832
rect 1797 2829 1821 2832
rect 1846 2829 1853 2832
rect 1857 2829 1879 2832
rect 1540 2819 1547 2822
rect 1551 2823 1570 2826
rect 1570 2816 1573 2822
rect 1598 2819 1605 2822
rect 1609 2823 1624 2826
rect 1672 2819 1679 2822
rect 1683 2823 1702 2826
rect 1702 2816 1705 2822
rect 1730 2819 1737 2822
rect 1741 2823 1756 2826
rect 1804 2819 1811 2822
rect 1815 2823 1834 2826
rect 1834 2816 1837 2822
rect 1862 2819 1869 2822
rect 1873 2823 1890 2826
rect 2469 2829 2474 2832
rect 2478 2829 2502 2832
rect 2527 2829 2534 2832
rect 2538 2829 2560 2832
rect 2580 2829 2587 2832
rect 2601 2829 2606 2832
rect 2610 2829 2634 2832
rect 2659 2829 2666 2832
rect 2670 2829 2692 2832
rect 2712 2829 2719 2832
rect 2733 2829 2738 2832
rect 2742 2829 2766 2832
rect 2791 2829 2798 2832
rect 2802 2829 2824 2832
rect 2485 2819 2492 2822
rect 2496 2823 2515 2826
rect 2515 2816 2518 2822
rect 2543 2819 2550 2822
rect 2554 2823 2569 2826
rect 2617 2819 2624 2822
rect 2628 2823 2647 2826
rect 2647 2816 2650 2822
rect 2675 2819 2682 2822
rect 2686 2823 2701 2826
rect 2749 2819 2756 2822
rect 2760 2823 2779 2826
rect 2779 2816 2782 2822
rect 2807 2819 2814 2822
rect 2818 2823 2835 2826
rect 1507 2800 1510 2812
rect 1528 2800 1531 2812
rect 1544 2800 1547 2812
rect 1558 2803 1570 2806
rect 1586 2800 1589 2812
rect 1602 2800 1605 2812
rect 1623 2800 1626 2812
rect 1639 2800 1642 2812
rect 1660 2800 1663 2812
rect 1676 2800 1679 2812
rect 1690 2803 1702 2806
rect 1718 2800 1721 2812
rect 1734 2800 1737 2812
rect 1755 2800 1758 2812
rect 1771 2800 1774 2812
rect 1792 2800 1795 2812
rect 1808 2800 1811 2812
rect 1822 2803 1834 2806
rect 1850 2800 1853 2812
rect 1866 2800 1869 2812
rect 1887 2800 1890 2812
rect 2452 2800 2455 2812
rect 2473 2800 2476 2812
rect 2489 2800 2492 2812
rect 2503 2803 2515 2806
rect 2531 2800 2534 2812
rect 2547 2800 2550 2812
rect 2568 2800 2571 2812
rect 2584 2800 2587 2812
rect 2605 2800 2608 2812
rect 2621 2800 2624 2812
rect 2635 2803 2647 2806
rect 2663 2800 2666 2812
rect 2679 2800 2682 2812
rect 2700 2800 2703 2812
rect 2716 2800 2719 2812
rect 2737 2800 2740 2812
rect 2753 2800 2756 2812
rect 2767 2803 2779 2806
rect 2795 2800 2798 2812
rect 2811 2800 2814 2812
rect 2832 2800 2835 2812
rect 1504 2796 1537 2800
rect 1541 2796 1565 2800
rect 1569 2796 1595 2800
rect 1599 2796 1669 2800
rect 1673 2796 1697 2800
rect 1701 2796 1727 2800
rect 1731 2796 1801 2800
rect 1805 2796 1829 2800
rect 1833 2796 1859 2800
rect 1863 2796 1916 2800
rect 2449 2796 2482 2800
rect 2486 2796 2510 2800
rect 2514 2796 2540 2800
rect 2544 2796 2614 2800
rect 2618 2796 2642 2800
rect 2646 2796 2672 2800
rect 2676 2796 2746 2800
rect 2750 2796 2774 2800
rect 2778 2796 2804 2800
rect 2808 2796 2861 2800
rect 1504 2789 1513 2793
rect 1517 2789 1564 2793
rect 1568 2789 1614 2793
rect 1618 2789 1645 2793
rect 1649 2789 1696 2793
rect 1700 2789 1746 2793
rect 1750 2789 1777 2793
rect 1781 2789 1828 2793
rect 1832 2789 1878 2793
rect 1882 2789 1952 2793
rect 2449 2789 2458 2793
rect 2462 2789 2509 2793
rect 2513 2789 2559 2793
rect 2563 2789 2590 2793
rect 2594 2789 2641 2793
rect 2645 2789 2691 2793
rect 2695 2789 2722 2793
rect 2726 2789 2773 2793
rect 2777 2789 2823 2793
rect 2827 2789 2897 2793
rect 1970 2781 1997 2785
rect 2001 2781 2033 2785
rect 2037 2781 2100 2785
rect 2104 2781 2129 2785
rect 2133 2781 2165 2785
rect 2169 2781 2232 2785
rect 2236 2781 2261 2785
rect 2265 2781 2297 2785
rect 2301 2781 2364 2785
rect 2368 2781 2393 2785
rect 2397 2781 2429 2785
rect 2433 2781 2496 2785
rect 2500 2781 2516 2785
rect 2915 2781 2942 2785
rect 2946 2781 2978 2785
rect 2982 2781 3045 2785
rect 3049 2781 3074 2785
rect 3078 2781 3110 2785
rect 3114 2781 3177 2785
rect 3181 2781 3206 2785
rect 3210 2781 3242 2785
rect 3246 2781 3309 2785
rect 3313 2781 3338 2785
rect 3342 2781 3374 2785
rect 3378 2781 3441 2785
rect 3445 2781 3461 2785
rect 1910 2774 2021 2778
rect 2025 2774 2049 2778
rect 2053 2774 2079 2778
rect 2083 2774 2116 2778
rect 2120 2774 2153 2778
rect 2157 2774 2181 2778
rect 2185 2774 2211 2778
rect 2215 2774 2248 2778
rect 2252 2774 2285 2778
rect 2289 2774 2313 2778
rect 2317 2774 2343 2778
rect 2347 2774 2380 2778
rect 2384 2774 2417 2778
rect 2421 2774 2445 2778
rect 2449 2774 2475 2778
rect 2479 2774 2512 2778
rect 2855 2774 2966 2778
rect 2970 2774 2994 2778
rect 2998 2774 3024 2778
rect 3028 2774 3061 2778
rect 3065 2774 3098 2778
rect 3102 2774 3126 2778
rect 3130 2774 3156 2778
rect 3160 2774 3193 2778
rect 3197 2774 3230 2778
rect 3234 2774 3258 2778
rect 3262 2774 3288 2778
rect 3292 2774 3325 2778
rect 3329 2774 3362 2778
rect 3366 2774 3390 2778
rect 3394 2774 3420 2778
rect 3424 2774 3457 2778
rect 1991 2764 1994 2774
rect 2012 2764 2015 2774
rect 2028 2764 2031 2774
rect 2042 2767 2047 2771
rect 2051 2767 2058 2771
rect 2070 2764 2073 2774
rect 2086 2764 2089 2774
rect 2107 2764 2110 2774
rect 2123 2764 2126 2774
rect 2144 2764 2147 2774
rect 2160 2764 2163 2774
rect 2174 2767 2179 2771
rect 2183 2767 2190 2771
rect 2202 2764 2205 2774
rect 2218 2764 2221 2774
rect 2239 2764 2242 2774
rect 2255 2764 2258 2774
rect 2276 2764 2279 2774
rect 2292 2764 2295 2774
rect 2306 2767 2311 2771
rect 2315 2767 2322 2771
rect 2334 2764 2337 2774
rect 2350 2764 2353 2774
rect 2371 2764 2374 2774
rect 2387 2764 2390 2774
rect 2408 2764 2411 2774
rect 2424 2764 2427 2774
rect 2438 2767 2443 2771
rect 2447 2767 2454 2771
rect 2466 2764 2469 2774
rect 2482 2764 2485 2774
rect 2503 2764 2506 2774
rect 2936 2764 2939 2774
rect 2957 2764 2960 2774
rect 2973 2764 2976 2774
rect 2987 2767 2992 2771
rect 2996 2767 3003 2771
rect 3015 2764 3018 2774
rect 3031 2764 3034 2774
rect 3052 2764 3055 2774
rect 3068 2764 3071 2774
rect 3089 2764 3092 2774
rect 3105 2764 3108 2774
rect 3119 2767 3124 2771
rect 3128 2767 3135 2771
rect 3147 2764 3150 2774
rect 3163 2764 3166 2774
rect 3184 2764 3187 2774
rect 3200 2764 3203 2774
rect 3221 2764 3224 2774
rect 3237 2764 3240 2774
rect 3251 2767 3256 2771
rect 3260 2767 3267 2771
rect 3279 2764 3282 2774
rect 3295 2764 3298 2774
rect 3316 2764 3319 2774
rect 3332 2764 3335 2774
rect 3353 2764 3356 2774
rect 3369 2764 3372 2774
rect 3383 2767 3388 2771
rect 3392 2767 3399 2771
rect 3411 2764 3414 2774
rect 3427 2764 3430 2774
rect 3448 2764 3451 2774
rect 1636 2748 1645 2752
rect 1649 2748 1681 2752
rect 1685 2748 1748 2752
rect 1752 2748 1964 2752
rect 2008 2750 2013 2753
rect 2017 2750 2041 2753
rect 2066 2750 2073 2753
rect 2077 2750 2099 2753
rect 1636 2741 1669 2745
rect 1673 2741 1697 2745
rect 1701 2741 1727 2745
rect 1731 2741 1764 2745
rect 1768 2741 1904 2745
rect 1639 2731 1642 2741
rect 1660 2731 1663 2741
rect 1676 2731 1679 2741
rect 1690 2734 1695 2738
rect 1699 2734 1706 2738
rect 1718 2731 1721 2741
rect 1734 2731 1737 2741
rect 1755 2731 1758 2741
rect 2024 2740 2031 2743
rect 2035 2744 2054 2747
rect 2054 2737 2057 2743
rect 2082 2740 2089 2743
rect 2093 2744 2110 2747
rect 2140 2750 2145 2753
rect 2149 2750 2173 2753
rect 2198 2750 2205 2753
rect 2209 2750 2231 2753
rect 2156 2740 2163 2743
rect 2167 2744 2186 2747
rect 2186 2737 2189 2743
rect 2214 2740 2221 2743
rect 2225 2744 2242 2747
rect 2272 2750 2277 2753
rect 2281 2750 2305 2753
rect 2330 2750 2337 2753
rect 2341 2750 2363 2753
rect 2288 2740 2295 2743
rect 2299 2744 2318 2747
rect 2318 2737 2321 2743
rect 2346 2740 2353 2743
rect 2357 2744 2374 2747
rect 2404 2750 2409 2753
rect 2413 2750 2437 2753
rect 2462 2750 2469 2753
rect 2473 2750 2495 2753
rect 2581 2748 2590 2752
rect 2594 2748 2626 2752
rect 2630 2748 2693 2752
rect 2697 2748 2909 2752
rect 2420 2740 2427 2743
rect 2431 2744 2450 2747
rect 1634 2714 1643 2718
rect 1656 2717 1661 2720
rect 1665 2717 1689 2720
rect 1714 2717 1721 2720
rect 1725 2717 1747 2720
rect 1991 2721 1994 2733
rect 2012 2721 2015 2733
rect 2028 2721 2031 2733
rect 2042 2724 2054 2727
rect 2070 2721 2073 2733
rect 2086 2721 2089 2733
rect 2107 2721 2110 2733
rect 2123 2721 2126 2733
rect 2144 2721 2147 2733
rect 2160 2721 2163 2733
rect 2174 2724 2186 2727
rect 2202 2721 2205 2733
rect 2218 2721 2221 2733
rect 2239 2721 2242 2733
rect 2255 2721 2258 2733
rect 2276 2721 2279 2733
rect 2292 2721 2295 2733
rect 2306 2724 2318 2727
rect 2334 2721 2337 2733
rect 2350 2721 2353 2733
rect 2371 2721 2374 2733
rect 2450 2737 2453 2743
rect 2478 2740 2485 2743
rect 2489 2744 2506 2747
rect 2953 2750 2958 2753
rect 2962 2750 2986 2753
rect 3011 2750 3018 2753
rect 3022 2750 3044 2753
rect 2581 2741 2614 2745
rect 2618 2741 2642 2745
rect 2646 2741 2672 2745
rect 2676 2741 2709 2745
rect 2713 2741 2849 2745
rect 2387 2721 2390 2733
rect 2408 2721 2411 2733
rect 2424 2721 2427 2733
rect 2438 2724 2450 2727
rect 2466 2721 2469 2733
rect 2482 2721 2485 2733
rect 2503 2721 2506 2733
rect 2584 2731 2587 2741
rect 2605 2731 2608 2741
rect 2621 2731 2624 2741
rect 2635 2734 2640 2738
rect 2644 2734 2651 2738
rect 2663 2731 2666 2741
rect 2679 2731 2682 2741
rect 2700 2731 2703 2741
rect 2969 2740 2976 2743
rect 2980 2744 2999 2747
rect 2999 2737 3002 2743
rect 3027 2740 3034 2743
rect 3038 2744 3055 2747
rect 3085 2750 3090 2753
rect 3094 2750 3118 2753
rect 3143 2750 3150 2753
rect 3154 2750 3176 2753
rect 3101 2740 3108 2743
rect 3112 2744 3131 2747
rect 3131 2737 3134 2743
rect 3159 2740 3166 2743
rect 3170 2744 3187 2747
rect 3217 2750 3222 2753
rect 3226 2750 3250 2753
rect 3275 2750 3282 2753
rect 3286 2750 3308 2753
rect 3233 2740 3240 2743
rect 3244 2744 3263 2747
rect 3263 2737 3266 2743
rect 3291 2740 3298 2743
rect 3302 2744 3319 2747
rect 3349 2750 3354 2753
rect 3358 2750 3382 2753
rect 3407 2750 3414 2753
rect 3418 2750 3440 2753
rect 3365 2740 3372 2743
rect 3376 2744 3395 2747
rect 1922 2717 2021 2721
rect 2025 2717 2049 2721
rect 2053 2717 2079 2721
rect 2083 2717 2153 2721
rect 2157 2717 2181 2721
rect 2185 2717 2211 2721
rect 2215 2717 2285 2721
rect 2289 2717 2313 2721
rect 2317 2717 2343 2721
rect 2347 2717 2417 2721
rect 2421 2717 2445 2721
rect 2449 2717 2475 2721
rect 2479 2717 2516 2721
rect 1672 2707 1679 2710
rect 1683 2711 1702 2714
rect 1702 2704 1705 2710
rect 1730 2707 1737 2710
rect 1741 2711 1756 2714
rect 2579 2714 2588 2718
rect 2601 2717 2606 2720
rect 2610 2717 2634 2720
rect 2659 2717 2666 2720
rect 2670 2717 2692 2720
rect 2936 2721 2939 2733
rect 2957 2721 2960 2733
rect 2973 2721 2976 2733
rect 2987 2724 2999 2727
rect 3015 2721 3018 2733
rect 3031 2721 3034 2733
rect 3052 2721 3055 2733
rect 3068 2721 3071 2733
rect 3089 2721 3092 2733
rect 3105 2721 3108 2733
rect 3119 2724 3131 2727
rect 3147 2721 3150 2733
rect 3163 2721 3166 2733
rect 3184 2721 3187 2733
rect 3200 2721 3203 2733
rect 3221 2721 3224 2733
rect 3237 2721 3240 2733
rect 3251 2724 3263 2727
rect 3279 2721 3282 2733
rect 3295 2721 3298 2733
rect 3316 2721 3319 2733
rect 3395 2737 3398 2743
rect 3423 2740 3430 2743
rect 3434 2744 3451 2747
rect 3332 2721 3335 2733
rect 3353 2721 3356 2733
rect 3369 2721 3372 2733
rect 3383 2724 3395 2727
rect 3411 2721 3414 2733
rect 3427 2721 3430 2733
rect 3448 2721 3451 2733
rect 2867 2717 2966 2721
rect 2970 2717 2994 2721
rect 2998 2717 3024 2721
rect 3028 2717 3098 2721
rect 3102 2717 3126 2721
rect 3130 2717 3156 2721
rect 3160 2717 3230 2721
rect 3234 2717 3258 2721
rect 3262 2717 3288 2721
rect 3292 2717 3362 2721
rect 3366 2717 3390 2721
rect 3394 2717 3420 2721
rect 3424 2717 3461 2721
rect 1958 2710 1997 2714
rect 2001 2710 2048 2714
rect 2052 2710 2098 2714
rect 2102 2710 2129 2714
rect 2133 2710 2180 2714
rect 2184 2710 2230 2714
rect 2234 2710 2261 2714
rect 2265 2710 2312 2714
rect 2316 2710 2362 2714
rect 2366 2710 2393 2714
rect 2397 2710 2444 2714
rect 2448 2710 2494 2714
rect 2498 2710 2516 2714
rect 2617 2707 2624 2710
rect 2628 2711 2647 2714
rect 1639 2688 1642 2700
rect 1660 2688 1663 2700
rect 1676 2688 1679 2700
rect 1690 2691 1702 2694
rect 1718 2688 1721 2700
rect 1734 2688 1737 2700
rect 1755 2688 1758 2700
rect 1910 2697 1995 2701
rect 1999 2697 2011 2701
rect 2015 2697 2029 2701
rect 2033 2697 2040 2701
rect 2044 2697 2046 2701
rect 2050 2697 2065 2701
rect 2069 2697 2102 2701
rect 2106 2697 2107 2701
rect 2111 2697 2119 2701
rect 2123 2697 2147 2701
rect 2151 2697 2163 2701
rect 2167 2697 2187 2701
rect 2191 2697 2241 2701
rect 2245 2697 2268 2701
rect 2272 2697 2322 2701
rect 2326 2697 2345 2701
rect 2647 2704 2650 2710
rect 2675 2707 2682 2710
rect 2686 2711 2701 2714
rect 2903 2710 2942 2714
rect 2946 2710 2993 2714
rect 2997 2710 3043 2714
rect 3047 2710 3074 2714
rect 3078 2710 3125 2714
rect 3129 2710 3175 2714
rect 3179 2710 3206 2714
rect 3210 2710 3257 2714
rect 3261 2710 3307 2714
rect 3311 2710 3338 2714
rect 3342 2710 3389 2714
rect 3393 2710 3439 2714
rect 3443 2710 3461 2714
rect 1946 2690 2022 2694
rect 2026 2690 2053 2694
rect 2057 2690 2075 2694
rect 2079 2690 2140 2694
rect 2144 2690 2158 2694
rect 2170 2693 2173 2697
rect 1636 2684 1669 2688
rect 1673 2684 1697 2688
rect 1701 2684 1727 2688
rect 1731 2684 1916 2688
rect 1636 2677 1645 2681
rect 1649 2677 1696 2681
rect 1700 2677 1746 2681
rect 1750 2677 1952 2681
rect 2065 2683 2068 2687
rect 2092 2683 2093 2687
rect 2137 2683 2139 2687
rect 2179 2680 2182 2685
rect 2194 2687 2197 2697
rect 2224 2693 2227 2697
rect 2251 2693 2254 2697
rect 1634 2661 1650 2665
rect 1759 2663 1763 2667
rect 1775 2663 1779 2667
rect 1783 2663 1989 2667
rect 1993 2663 1997 2667
rect 2005 2666 2008 2672
rect 2012 2666 2015 2672
rect 2005 2663 2015 2666
rect 2005 2658 2008 2663
rect 1642 2654 1646 2658
rect 1658 2654 1779 2658
rect 2012 2658 2015 2663
rect 2021 2668 2024 2672
rect 2021 2664 2023 2668
rect 2027 2664 2029 2668
rect 2037 2667 2040 2672
rect 2065 2669 2068 2672
rect 2037 2665 2048 2667
rect 2021 2658 2024 2664
rect 2037 2663 2043 2665
rect 2037 2658 2040 2663
rect 2047 2663 2048 2665
rect 2066 2665 2068 2669
rect 2065 2658 2068 2665
rect 2168 2676 2171 2679
rect 2210 2676 2213 2679
rect 2081 2668 2084 2672
rect 2091 2668 2094 2672
rect 2091 2664 2100 2668
rect 2112 2667 2115 2672
rect 2137 2668 2140 2672
rect 2081 2658 2084 2664
rect 2091 2658 2094 2664
rect 2112 2663 2113 2667
rect 2117 2663 2120 2666
rect 2139 2664 2140 2668
rect 2155 2667 2158 2672
rect 2179 2671 2182 2676
rect 2187 2672 2198 2675
rect 2210 2673 2218 2676
rect 2112 2658 2115 2663
rect 2137 2658 2140 2664
rect 2155 2658 2158 2663
rect 1629 2646 1645 2650
rect 1649 2646 1712 2650
rect 1716 2646 1748 2650
rect 1752 2646 1964 2650
rect 2057 2645 2058 2649
rect 2082 2646 2083 2650
rect 2129 2645 2130 2649
rect 1633 2639 1666 2643
rect 1670 2639 1696 2643
rect 1700 2639 1724 2643
rect 1728 2639 1904 2643
rect 1639 2629 1642 2639
rect 1660 2629 1663 2639
rect 1676 2629 1679 2639
rect 1691 2632 1698 2636
rect 1702 2632 1707 2636
rect 1718 2629 1721 2639
rect 1734 2629 1737 2639
rect 1755 2629 1758 2639
rect 1934 2638 2010 2642
rect 2014 2638 2069 2642
rect 2073 2638 2094 2642
rect 2098 2638 2125 2642
rect 2129 2638 2158 2642
rect 2170 2635 2173 2667
rect 2187 2666 2190 2672
rect 2210 2667 2213 2673
rect 2222 2668 2225 2671
rect 2233 2671 2236 2685
rect 2260 2680 2263 2685
rect 2275 2687 2278 2697
rect 2305 2693 2308 2697
rect 2244 2676 2245 2679
rect 2249 2676 2252 2679
rect 2584 2688 2587 2700
rect 2605 2688 2608 2700
rect 2621 2688 2624 2700
rect 2635 2691 2647 2694
rect 2663 2688 2666 2700
rect 2679 2688 2682 2700
rect 2700 2688 2703 2700
rect 2855 2697 2940 2701
rect 2944 2697 2956 2701
rect 2960 2697 2974 2701
rect 2978 2697 2985 2701
rect 2989 2697 2991 2701
rect 2995 2697 3010 2701
rect 3014 2697 3047 2701
rect 3051 2697 3052 2701
rect 3056 2697 3064 2701
rect 3068 2697 3092 2701
rect 3096 2697 3108 2701
rect 3112 2697 3132 2701
rect 3136 2697 3186 2701
rect 3190 2697 3213 2701
rect 3217 2697 3267 2701
rect 3271 2697 3290 2701
rect 2891 2690 2967 2694
rect 2971 2690 2998 2694
rect 3002 2690 3020 2694
rect 3024 2690 3085 2694
rect 3089 2690 3103 2694
rect 3115 2693 3118 2697
rect 2291 2676 2294 2679
rect 2233 2668 2241 2671
rect 2260 2671 2263 2676
rect 2233 2663 2236 2668
rect 2241 2664 2245 2668
rect 2268 2672 2279 2675
rect 2291 2673 2299 2676
rect 2185 2657 2190 2662
rect 2194 2635 2197 2663
rect 2224 2635 2227 2659
rect 2251 2635 2254 2667
rect 2268 2666 2271 2672
rect 2291 2667 2294 2673
rect 2303 2668 2306 2671
rect 2314 2671 2317 2685
rect 2581 2684 2614 2688
rect 2618 2684 2642 2688
rect 2646 2684 2672 2688
rect 2676 2684 2861 2688
rect 2581 2677 2590 2681
rect 2594 2677 2641 2681
rect 2645 2677 2691 2681
rect 2695 2677 2897 2681
rect 3010 2683 3013 2687
rect 3037 2683 3038 2687
rect 3082 2683 3084 2687
rect 3124 2680 3127 2685
rect 3139 2687 3142 2697
rect 3169 2693 3172 2697
rect 3196 2693 3199 2697
rect 2314 2668 2326 2671
rect 2314 2663 2317 2668
rect 2266 2657 2271 2662
rect 2275 2635 2278 2663
rect 2579 2661 2595 2665
rect 2704 2663 2708 2667
rect 2720 2663 2724 2667
rect 2728 2663 2934 2667
rect 2938 2663 2942 2667
rect 2950 2666 2953 2672
rect 2957 2666 2960 2672
rect 2950 2663 2960 2666
rect 2305 2635 2308 2659
rect 2950 2658 2953 2663
rect 2587 2654 2591 2658
rect 2603 2654 2724 2658
rect 2957 2658 2960 2663
rect 2966 2668 2969 2672
rect 2966 2664 2968 2668
rect 2972 2664 2974 2668
rect 2982 2667 2985 2672
rect 3010 2669 3013 2672
rect 2982 2665 2993 2667
rect 2966 2658 2969 2664
rect 2982 2663 2988 2665
rect 2982 2658 2985 2663
rect 2992 2663 2993 2665
rect 3011 2665 3013 2669
rect 3010 2658 3013 2665
rect 3113 2676 3116 2679
rect 3155 2676 3158 2679
rect 3026 2668 3029 2672
rect 3036 2668 3039 2672
rect 3036 2664 3045 2668
rect 3057 2667 3060 2672
rect 3082 2668 3085 2672
rect 3026 2658 3029 2664
rect 3036 2658 3039 2664
rect 3057 2663 3058 2667
rect 3062 2663 3065 2666
rect 3084 2664 3085 2668
rect 3100 2667 3103 2672
rect 3124 2671 3127 2676
rect 3132 2672 3143 2675
rect 3155 2673 3163 2676
rect 3057 2658 3060 2663
rect 3082 2658 3085 2664
rect 3100 2658 3103 2663
rect 2574 2646 2590 2650
rect 2594 2646 2657 2650
rect 2661 2646 2693 2650
rect 2697 2646 2909 2650
rect 3002 2645 3003 2649
rect 3027 2646 3028 2650
rect 3074 2645 3075 2649
rect 2578 2639 2611 2643
rect 2615 2639 2641 2643
rect 2645 2639 2669 2643
rect 2673 2639 2849 2643
rect 1922 2631 1996 2635
rect 2000 2631 2002 2635
rect 2006 2631 2010 2635
rect 2014 2631 2028 2635
rect 2032 2631 2037 2635
rect 2041 2631 2046 2635
rect 2050 2631 2069 2635
rect 2073 2631 2103 2635
rect 2107 2631 2118 2635
rect 2122 2631 2146 2635
rect 2150 2631 2163 2635
rect 2167 2631 2187 2635
rect 2191 2631 2241 2635
rect 2248 2631 2268 2635
rect 2272 2631 2322 2635
rect 1650 2615 1672 2618
rect 1676 2615 1683 2618
rect 1934 2624 2010 2628
rect 2014 2624 2069 2628
rect 2073 2624 2094 2628
rect 2098 2624 2125 2628
rect 2129 2624 2158 2628
rect 1708 2615 1732 2618
rect 1736 2615 1741 2618
rect 2057 2617 2058 2621
rect 2082 2616 2083 2620
rect 2129 2617 2130 2621
rect 1754 2612 1763 2616
rect 1641 2609 1656 2612
rect 1695 2609 1714 2612
rect 1660 2605 1667 2608
rect 1692 2602 1695 2608
rect 1718 2605 1725 2608
rect 2005 2603 2008 2608
rect 2012 2603 2015 2608
rect 1995 2600 1997 2603
rect 2005 2600 2015 2603
rect 1639 2586 1642 2598
rect 1660 2586 1663 2598
rect 1676 2586 1679 2598
rect 1695 2589 1707 2592
rect 1718 2586 1721 2598
rect 1734 2586 1737 2598
rect 1755 2586 1758 2598
rect 2005 2594 2008 2600
rect 2012 2594 2015 2600
rect 2021 2602 2024 2608
rect 2037 2603 2040 2608
rect 2021 2598 2023 2602
rect 2027 2598 2029 2602
rect 2037 2601 2043 2603
rect 2047 2601 2048 2603
rect 2037 2599 2048 2601
rect 2065 2601 2068 2608
rect 2021 2594 2024 2598
rect 2037 2594 2040 2599
rect 2066 2597 2068 2601
rect 2065 2594 2068 2597
rect 2081 2602 2084 2608
rect 2091 2602 2094 2608
rect 2112 2603 2115 2608
rect 2091 2598 2100 2602
rect 2112 2599 2113 2603
rect 2117 2600 2120 2603
rect 2137 2602 2140 2608
rect 2155 2603 2158 2608
rect 2194 2611 2197 2631
rect 2275 2611 2278 2631
rect 2584 2629 2587 2639
rect 2605 2629 2608 2639
rect 2621 2629 2624 2639
rect 2636 2632 2643 2636
rect 2647 2632 2652 2636
rect 2663 2629 2666 2639
rect 2679 2629 2682 2639
rect 2700 2629 2703 2639
rect 2879 2638 2955 2642
rect 2959 2638 3014 2642
rect 3018 2638 3039 2642
rect 3043 2638 3070 2642
rect 3074 2638 3103 2642
rect 3115 2635 3118 2667
rect 3132 2666 3135 2672
rect 3155 2667 3158 2673
rect 3167 2668 3170 2671
rect 3178 2671 3181 2685
rect 3205 2680 3208 2685
rect 3220 2687 3223 2697
rect 3250 2693 3253 2697
rect 3189 2676 3190 2679
rect 3194 2676 3197 2679
rect 3236 2676 3239 2679
rect 3178 2668 3186 2671
rect 3205 2671 3208 2676
rect 3178 2663 3181 2668
rect 3186 2664 3190 2668
rect 3213 2672 3224 2675
rect 3236 2673 3244 2676
rect 3130 2657 3135 2662
rect 3139 2635 3142 2663
rect 3169 2635 3172 2659
rect 3196 2635 3199 2667
rect 3213 2666 3216 2672
rect 3236 2667 3239 2673
rect 3248 2668 3251 2671
rect 3259 2671 3262 2685
rect 3259 2668 3271 2671
rect 3259 2663 3262 2668
rect 3211 2657 3216 2662
rect 3220 2635 3223 2663
rect 3250 2635 3253 2659
rect 2867 2631 2941 2635
rect 2945 2631 2947 2635
rect 2951 2631 2955 2635
rect 2959 2631 2973 2635
rect 2977 2631 2982 2635
rect 2986 2631 2991 2635
rect 2995 2631 3014 2635
rect 3018 2631 3048 2635
rect 3052 2631 3063 2635
rect 3067 2631 3091 2635
rect 3095 2631 3108 2635
rect 3112 2631 3132 2635
rect 3136 2631 3186 2635
rect 3193 2631 3213 2635
rect 3217 2631 3267 2635
rect 2595 2615 2617 2618
rect 2621 2615 2628 2618
rect 2879 2624 2955 2628
rect 2959 2624 3014 2628
rect 3018 2624 3039 2628
rect 3043 2624 3070 2628
rect 3074 2624 3103 2628
rect 2653 2615 2677 2618
rect 2681 2615 2686 2618
rect 3002 2617 3003 2621
rect 3027 2616 3028 2620
rect 3074 2617 3075 2621
rect 2699 2612 2708 2616
rect 2586 2609 2601 2612
rect 2081 2594 2084 2598
rect 2091 2594 2094 2598
rect 2112 2594 2115 2599
rect 2139 2598 2140 2602
rect 2137 2594 2140 2598
rect 2155 2594 2158 2599
rect 2185 2598 2190 2603
rect 2194 2599 2195 2602
rect 2210 2601 2213 2607
rect 2210 2598 2218 2601
rect 2265 2598 2270 2603
rect 2274 2599 2276 2602
rect 2291 2601 2294 2607
rect 2640 2609 2659 2612
rect 2605 2605 2612 2608
rect 2637 2602 2640 2608
rect 2291 2598 2299 2601
rect 2663 2605 2670 2608
rect 2950 2603 2953 2608
rect 2957 2603 2960 2608
rect 2940 2600 2942 2603
rect 2950 2600 2960 2603
rect 2210 2595 2213 2598
rect 2291 2595 2294 2598
rect 1629 2582 1666 2586
rect 1670 2582 1696 2586
rect 1700 2582 1724 2586
rect 1728 2582 1916 2586
rect 2065 2579 2068 2583
rect 2092 2579 2093 2583
rect 2137 2579 2139 2583
rect 1629 2575 1647 2579
rect 1651 2575 1697 2579
rect 1701 2575 1748 2579
rect 1752 2575 1952 2579
rect 2010 2572 2022 2576
rect 2026 2572 2053 2576
rect 2057 2572 2075 2576
rect 2079 2572 2140 2576
rect 2144 2572 2158 2576
rect 2194 2569 2197 2587
rect 2275 2569 2278 2587
rect 2584 2586 2587 2598
rect 2605 2586 2608 2598
rect 2621 2586 2624 2598
rect 2640 2589 2652 2592
rect 2663 2586 2666 2598
rect 2679 2586 2682 2598
rect 2700 2586 2703 2598
rect 2950 2594 2953 2600
rect 2957 2594 2960 2600
rect 2966 2602 2969 2608
rect 2982 2603 2985 2608
rect 2966 2598 2968 2602
rect 2972 2598 2974 2602
rect 2982 2601 2988 2603
rect 2992 2601 2993 2603
rect 2982 2599 2993 2601
rect 3010 2601 3013 2608
rect 2966 2594 2969 2598
rect 2982 2594 2985 2599
rect 3011 2597 3013 2601
rect 3010 2594 3013 2597
rect 3026 2602 3029 2608
rect 3036 2602 3039 2608
rect 3057 2603 3060 2608
rect 3036 2598 3045 2602
rect 3057 2599 3058 2603
rect 3062 2600 3065 2603
rect 3082 2602 3085 2608
rect 3100 2603 3103 2608
rect 3139 2611 3142 2631
rect 3220 2611 3223 2631
rect 3026 2594 3029 2598
rect 3036 2594 3039 2598
rect 3057 2594 3060 2599
rect 3084 2598 3085 2602
rect 3082 2594 3085 2598
rect 3100 2594 3103 2599
rect 3130 2598 3135 2603
rect 3139 2599 3140 2602
rect 3155 2601 3158 2607
rect 3155 2598 3163 2601
rect 3210 2598 3215 2603
rect 3219 2599 3221 2602
rect 3236 2601 3239 2607
rect 3236 2598 3244 2601
rect 3155 2595 3158 2598
rect 3236 2595 3239 2598
rect 2574 2582 2611 2586
rect 2615 2582 2641 2586
rect 2645 2582 2669 2586
rect 2673 2582 2861 2586
rect 3010 2579 3013 2583
rect 3037 2579 3038 2583
rect 3082 2579 3084 2583
rect 2574 2575 2592 2579
rect 2596 2575 2642 2579
rect 2646 2575 2693 2579
rect 2697 2575 2897 2579
rect 2955 2572 2967 2576
rect 2971 2572 2998 2576
rect 3002 2572 3020 2576
rect 3024 2572 3085 2576
rect 3089 2572 3103 2576
rect 3139 2569 3142 2587
rect 3220 2569 3223 2587
rect 1910 2565 1995 2569
rect 1999 2565 2011 2569
rect 2015 2565 2029 2569
rect 2033 2565 2040 2569
rect 2044 2565 2046 2569
rect 2050 2565 2065 2569
rect 2069 2565 2102 2569
rect 2106 2565 2107 2569
rect 2111 2565 2119 2569
rect 2123 2565 2147 2569
rect 2151 2565 2163 2569
rect 2167 2565 2187 2569
rect 2191 2565 2241 2569
rect 2245 2565 2268 2569
rect 2272 2565 2330 2569
rect 2334 2565 2345 2569
rect 2855 2565 2940 2569
rect 2944 2565 2956 2569
rect 2960 2565 2974 2569
rect 2978 2565 2985 2569
rect 2989 2565 2991 2569
rect 2995 2565 3010 2569
rect 3014 2565 3047 2569
rect 3051 2565 3052 2569
rect 3056 2565 3064 2569
rect 3068 2565 3092 2569
rect 3096 2565 3108 2569
rect 3112 2565 3132 2569
rect 3136 2565 3186 2569
rect 3190 2565 3213 2569
rect 3217 2565 3275 2569
rect 3279 2565 3290 2569
rect 1946 2558 2006 2562
rect 2010 2558 2022 2562
rect 2026 2558 2053 2562
rect 2057 2558 2075 2562
rect 2079 2558 2140 2562
rect 2144 2558 2158 2562
rect 2194 2555 2197 2565
rect 2224 2561 2227 2565
rect 2275 2561 2278 2565
rect 2065 2551 2068 2555
rect 2092 2551 2093 2555
rect 2137 2551 2139 2555
rect 1994 2531 1997 2534
rect 2005 2534 2008 2540
rect 2012 2534 2015 2540
rect 2005 2531 2015 2534
rect 2005 2526 2008 2531
rect 2012 2526 2015 2531
rect 2021 2536 2024 2540
rect 2021 2532 2023 2536
rect 2027 2532 2029 2536
rect 2037 2535 2040 2540
rect 2065 2537 2068 2540
rect 2037 2533 2048 2535
rect 2021 2526 2024 2532
rect 2037 2531 2043 2533
rect 2037 2526 2040 2531
rect 2047 2531 2048 2533
rect 2066 2533 2068 2537
rect 2065 2526 2068 2533
rect 2210 2544 2213 2547
rect 2081 2536 2084 2540
rect 2091 2536 2094 2540
rect 2091 2532 2100 2536
rect 2112 2535 2115 2540
rect 2137 2536 2140 2540
rect 2081 2526 2084 2532
rect 2091 2526 2094 2532
rect 2112 2531 2113 2535
rect 2117 2531 2120 2534
rect 2139 2532 2140 2536
rect 2155 2535 2158 2540
rect 2187 2540 2198 2543
rect 2210 2541 2218 2544
rect 2112 2526 2115 2531
rect 2137 2526 2140 2532
rect 2187 2534 2190 2540
rect 2210 2535 2213 2541
rect 2222 2536 2225 2539
rect 2233 2539 2236 2553
rect 2284 2548 2287 2553
rect 2299 2555 2302 2565
rect 2329 2561 2332 2565
rect 2268 2544 2269 2547
rect 2273 2544 2276 2547
rect 2891 2558 2951 2562
rect 2955 2558 2967 2562
rect 2971 2558 2998 2562
rect 3002 2558 3020 2562
rect 3024 2558 3085 2562
rect 3089 2558 3103 2562
rect 3139 2555 3142 2565
rect 3169 2561 3172 2565
rect 3220 2561 3223 2565
rect 2315 2544 2318 2547
rect 2241 2539 2246 2544
rect 2284 2539 2287 2544
rect 2233 2536 2241 2539
rect 2155 2526 2158 2531
rect 2233 2531 2236 2536
rect 2292 2540 2303 2543
rect 2315 2541 2323 2544
rect 2185 2525 2190 2530
rect 2057 2513 2058 2517
rect 2082 2514 2083 2518
rect 2129 2513 2130 2517
rect 1934 2506 2010 2510
rect 2014 2506 2069 2510
rect 2073 2506 2094 2510
rect 2098 2506 2125 2510
rect 2129 2506 2158 2510
rect 2194 2503 2197 2531
rect 2224 2503 2227 2527
rect 2275 2503 2278 2535
rect 2292 2534 2295 2540
rect 2315 2535 2318 2541
rect 2327 2536 2330 2539
rect 2338 2539 2341 2553
rect 3010 2551 3013 2555
rect 3037 2551 3038 2555
rect 3082 2551 3084 2555
rect 2338 2536 2344 2539
rect 2338 2531 2341 2536
rect 2939 2531 2942 2534
rect 2950 2534 2953 2540
rect 2957 2534 2960 2540
rect 2950 2531 2960 2534
rect 2290 2525 2295 2530
rect 2299 2503 2302 2531
rect 2329 2503 2332 2527
rect 2950 2526 2953 2531
rect 2957 2526 2960 2531
rect 2966 2536 2969 2540
rect 2966 2532 2968 2536
rect 2972 2532 2974 2536
rect 2982 2535 2985 2540
rect 3010 2537 3013 2540
rect 2982 2533 2993 2535
rect 2966 2526 2969 2532
rect 2982 2531 2988 2533
rect 2982 2526 2985 2531
rect 2992 2531 2993 2533
rect 3011 2533 3013 2537
rect 3010 2526 3013 2533
rect 3155 2544 3158 2547
rect 3026 2536 3029 2540
rect 3036 2536 3039 2540
rect 3036 2532 3045 2536
rect 3057 2535 3060 2540
rect 3082 2536 3085 2540
rect 3026 2526 3029 2532
rect 3036 2526 3039 2532
rect 3057 2531 3058 2535
rect 3062 2531 3065 2534
rect 3084 2532 3085 2536
rect 3100 2535 3103 2540
rect 3132 2540 3143 2543
rect 3155 2541 3163 2544
rect 3057 2526 3060 2531
rect 3082 2526 3085 2532
rect 3132 2534 3135 2540
rect 3155 2535 3158 2541
rect 3167 2536 3170 2539
rect 3178 2539 3181 2553
rect 3229 2548 3232 2553
rect 3244 2555 3247 2565
rect 3274 2561 3277 2565
rect 3213 2544 3214 2547
rect 3218 2544 3221 2547
rect 3260 2544 3263 2547
rect 3186 2539 3191 2544
rect 3229 2539 3232 2544
rect 3178 2536 3186 2539
rect 3100 2526 3103 2531
rect 3178 2531 3181 2536
rect 3237 2540 3248 2543
rect 3260 2541 3268 2544
rect 3130 2525 3135 2530
rect 3002 2513 3003 2517
rect 3027 2514 3028 2518
rect 3074 2513 3075 2517
rect 2879 2506 2955 2510
rect 2959 2506 3014 2510
rect 3018 2506 3039 2510
rect 3043 2506 3070 2510
rect 3074 2506 3103 2510
rect 3139 2503 3142 2531
rect 3169 2503 3172 2527
rect 3220 2503 3223 2535
rect 3237 2534 3240 2540
rect 3260 2535 3263 2541
rect 3272 2536 3275 2539
rect 3283 2539 3286 2553
rect 3283 2536 3289 2539
rect 3283 2531 3286 2536
rect 3235 2525 3240 2530
rect 3244 2503 3247 2531
rect 3274 2503 3277 2527
rect 1922 2499 1996 2503
rect 2000 2499 2002 2503
rect 2006 2499 2010 2503
rect 2014 2499 2028 2503
rect 2032 2499 2037 2503
rect 2041 2499 2046 2503
rect 2050 2499 2069 2503
rect 2073 2499 2103 2503
rect 2107 2499 2118 2503
rect 2122 2499 2146 2503
rect 2150 2499 2163 2503
rect 2167 2499 2187 2503
rect 2191 2499 2241 2503
rect 2245 2499 2268 2503
rect 2272 2499 2292 2503
rect 2296 2499 2344 2503
rect 2867 2499 2941 2503
rect 2945 2499 2947 2503
rect 2951 2499 2955 2503
rect 2959 2499 2973 2503
rect 2977 2499 2982 2503
rect 2986 2499 2991 2503
rect 2995 2499 3014 2503
rect 3018 2499 3048 2503
rect 3052 2499 3063 2503
rect 3067 2499 3091 2503
rect 3095 2499 3108 2503
rect 3112 2499 3132 2503
rect 3136 2499 3186 2503
rect 3190 2499 3213 2503
rect 3217 2499 3237 2503
rect 3241 2499 3289 2503
rect 1934 2492 2010 2496
rect 2014 2492 2069 2496
rect 2073 2492 2094 2496
rect 2098 2492 2125 2496
rect 2129 2492 2158 2496
rect 2057 2485 2058 2489
rect 2082 2484 2083 2488
rect 2129 2485 2130 2489
rect 2194 2480 2197 2499
rect 2299 2480 2302 2499
rect 2879 2492 2955 2496
rect 2959 2492 3014 2496
rect 3018 2492 3039 2496
rect 3043 2492 3070 2496
rect 3074 2492 3103 2496
rect 3002 2485 3003 2489
rect 3027 2484 3028 2488
rect 3074 2485 3075 2489
rect 3139 2480 3142 2499
rect 3244 2480 3247 2499
rect 2005 2471 2008 2476
rect 2012 2471 2015 2476
rect 1995 2468 1997 2471
rect 2005 2468 2015 2471
rect 2005 2462 2008 2468
rect 2012 2462 2015 2468
rect 2021 2470 2024 2476
rect 2037 2471 2040 2476
rect 2021 2466 2023 2470
rect 2027 2466 2029 2470
rect 2037 2469 2043 2471
rect 2047 2469 2048 2471
rect 2037 2467 2048 2469
rect 2065 2469 2068 2476
rect 2021 2462 2024 2466
rect 2037 2462 2040 2467
rect 2066 2465 2068 2469
rect 2065 2462 2068 2465
rect 2081 2470 2084 2476
rect 2091 2470 2094 2476
rect 2112 2471 2115 2476
rect 2091 2466 2100 2470
rect 2112 2467 2113 2471
rect 2117 2468 2120 2471
rect 2137 2470 2140 2476
rect 2155 2471 2158 2476
rect 2081 2462 2084 2466
rect 2091 2462 2094 2466
rect 2112 2462 2115 2467
rect 2139 2466 2140 2470
rect 2184 2467 2189 2472
rect 2193 2468 2195 2471
rect 2210 2470 2213 2476
rect 2210 2467 2218 2470
rect 2290 2467 2295 2472
rect 2299 2468 2300 2471
rect 2315 2470 2318 2476
rect 2315 2467 2323 2470
rect 2950 2471 2953 2476
rect 2957 2471 2960 2476
rect 2940 2468 2942 2471
rect 2950 2468 2960 2471
rect 2137 2462 2140 2466
rect 2155 2462 2158 2467
rect 2210 2464 2213 2467
rect 2315 2464 2318 2467
rect 2950 2462 2953 2468
rect 2065 2447 2068 2451
rect 2092 2447 2093 2451
rect 2137 2447 2139 2451
rect 1946 2440 2022 2444
rect 2026 2440 2053 2444
rect 2057 2440 2075 2444
rect 2079 2440 2140 2444
rect 2144 2440 2158 2444
rect 2194 2437 2197 2456
rect 2299 2437 2302 2456
rect 2957 2462 2960 2468
rect 2966 2470 2969 2476
rect 2982 2471 2985 2476
rect 2966 2466 2968 2470
rect 2972 2466 2974 2470
rect 2982 2469 2988 2471
rect 2992 2469 2993 2471
rect 2982 2467 2993 2469
rect 3010 2469 3013 2476
rect 2966 2462 2969 2466
rect 2982 2462 2985 2467
rect 3011 2465 3013 2469
rect 3010 2462 3013 2465
rect 3026 2470 3029 2476
rect 3036 2470 3039 2476
rect 3057 2471 3060 2476
rect 3036 2466 3045 2470
rect 3057 2467 3058 2471
rect 3062 2468 3065 2471
rect 3082 2470 3085 2476
rect 3100 2471 3103 2476
rect 3026 2462 3029 2466
rect 3036 2462 3039 2466
rect 3057 2462 3060 2467
rect 3084 2466 3085 2470
rect 3129 2467 3134 2472
rect 3138 2468 3140 2471
rect 3155 2470 3158 2476
rect 3155 2467 3163 2470
rect 3235 2467 3240 2472
rect 3244 2468 3245 2471
rect 3260 2470 3263 2476
rect 3260 2467 3268 2470
rect 3082 2462 3085 2466
rect 3100 2462 3103 2467
rect 3155 2464 3158 2467
rect 3260 2464 3263 2467
rect 3010 2447 3013 2451
rect 3037 2447 3038 2451
rect 3082 2447 3084 2451
rect 2891 2440 2967 2444
rect 2971 2440 2998 2444
rect 3002 2440 3020 2444
rect 3024 2440 3085 2444
rect 3089 2440 3103 2444
rect 3139 2437 3142 2456
rect 3244 2437 3247 2456
rect 1910 2433 1995 2437
rect 1999 2433 2011 2437
rect 2015 2433 2029 2437
rect 2033 2433 2040 2437
rect 2044 2433 2046 2437
rect 2050 2433 2065 2437
rect 2069 2433 2102 2437
rect 2106 2433 2107 2437
rect 2111 2433 2119 2437
rect 2123 2433 2147 2437
rect 2151 2433 2163 2437
rect 2167 2433 2187 2437
rect 2191 2433 2241 2437
rect 2245 2433 2268 2437
rect 2272 2433 2322 2437
rect 2326 2433 2330 2437
rect 2334 2433 2358 2437
rect 2362 2433 2412 2437
rect 2855 2433 2940 2437
rect 2944 2433 2956 2437
rect 2960 2433 2974 2437
rect 2978 2433 2985 2437
rect 2989 2433 2991 2437
rect 2995 2433 3010 2437
rect 3014 2433 3047 2437
rect 3051 2433 3052 2437
rect 3056 2433 3064 2437
rect 3068 2433 3092 2437
rect 3096 2433 3108 2437
rect 3112 2433 3132 2437
rect 3136 2433 3186 2437
rect 3190 2433 3213 2437
rect 3217 2433 3267 2437
rect 3271 2433 3275 2437
rect 3279 2433 3303 2437
rect 3307 2433 3357 2437
rect 1946 2426 2022 2430
rect 2026 2426 2053 2430
rect 2057 2426 2075 2430
rect 2079 2426 2140 2430
rect 2144 2426 2158 2430
rect 2194 2423 2197 2433
rect 2224 2429 2227 2433
rect 2251 2429 2254 2433
rect 2065 2419 2068 2423
rect 2092 2419 2093 2423
rect 2137 2419 2139 2423
rect 1994 2399 1997 2402
rect 2005 2402 2008 2408
rect 2012 2402 2015 2408
rect 2005 2399 2015 2402
rect 2005 2394 2008 2399
rect 2012 2394 2015 2399
rect 2021 2404 2024 2408
rect 2021 2400 2023 2404
rect 2027 2400 2029 2404
rect 2037 2403 2040 2408
rect 2065 2405 2068 2408
rect 2037 2401 2048 2403
rect 2021 2394 2024 2400
rect 2037 2399 2043 2401
rect 2037 2394 2040 2399
rect 2047 2399 2048 2401
rect 2066 2401 2068 2405
rect 2065 2394 2068 2401
rect 2210 2412 2213 2415
rect 2081 2404 2084 2408
rect 2091 2404 2094 2408
rect 2091 2400 2100 2404
rect 2112 2403 2115 2408
rect 2137 2404 2140 2408
rect 2081 2394 2084 2400
rect 2091 2394 2094 2400
rect 2112 2399 2113 2403
rect 2117 2399 2120 2402
rect 2139 2400 2140 2404
rect 2155 2403 2158 2408
rect 2187 2408 2198 2411
rect 2210 2409 2218 2412
rect 2112 2394 2115 2399
rect 2137 2394 2140 2400
rect 2187 2402 2190 2408
rect 2210 2403 2213 2409
rect 2222 2404 2225 2407
rect 2233 2407 2236 2421
rect 2260 2416 2263 2421
rect 2275 2423 2278 2433
rect 2305 2429 2308 2433
rect 2341 2429 2344 2433
rect 2244 2412 2245 2415
rect 2249 2412 2252 2415
rect 2291 2412 2294 2415
rect 2233 2404 2241 2407
rect 2260 2407 2263 2412
rect 2155 2394 2158 2399
rect 2233 2399 2236 2404
rect 2241 2400 2245 2404
rect 2268 2408 2279 2411
rect 2291 2409 2299 2412
rect 2185 2393 2190 2398
rect 2057 2381 2058 2385
rect 2082 2382 2083 2386
rect 2129 2381 2130 2385
rect 1934 2374 2010 2378
rect 2014 2374 2069 2378
rect 2073 2374 2094 2378
rect 2098 2374 2125 2378
rect 2129 2374 2158 2378
rect 2194 2371 2197 2399
rect 2224 2371 2227 2395
rect 2251 2371 2254 2403
rect 2268 2402 2271 2408
rect 2291 2403 2294 2409
rect 2303 2404 2306 2407
rect 2314 2407 2317 2421
rect 2350 2416 2353 2421
rect 2365 2423 2368 2433
rect 2395 2429 2398 2433
rect 2339 2412 2342 2415
rect 2891 2426 2967 2430
rect 2971 2426 2998 2430
rect 3002 2426 3020 2430
rect 3024 2426 3085 2430
rect 3089 2426 3103 2430
rect 3139 2423 3142 2433
rect 3169 2429 3172 2433
rect 3196 2429 3199 2433
rect 2381 2412 2384 2415
rect 2314 2404 2323 2407
rect 2350 2407 2353 2412
rect 2314 2399 2317 2404
rect 2266 2393 2271 2398
rect 2275 2371 2278 2399
rect 2357 2410 2369 2411
rect 2361 2408 2369 2410
rect 2381 2409 2389 2412
rect 2381 2403 2384 2409
rect 2393 2404 2396 2407
rect 2404 2407 2407 2421
rect 3010 2419 3013 2423
rect 3037 2419 3038 2423
rect 3082 2419 3084 2423
rect 2404 2404 2424 2407
rect 2305 2371 2308 2395
rect 2341 2371 2344 2403
rect 2404 2399 2407 2404
rect 2939 2399 2942 2402
rect 2950 2402 2953 2408
rect 2957 2402 2960 2408
rect 2950 2399 2960 2402
rect 2365 2371 2368 2399
rect 2395 2371 2398 2395
rect 2950 2394 2953 2399
rect 2957 2394 2960 2399
rect 2966 2404 2969 2408
rect 2966 2400 2968 2404
rect 2972 2400 2974 2404
rect 2982 2403 2985 2408
rect 3010 2405 3013 2408
rect 2982 2401 2993 2403
rect 2966 2394 2969 2400
rect 2982 2399 2988 2401
rect 2982 2394 2985 2399
rect 2992 2399 2993 2401
rect 3011 2401 3013 2405
rect 3010 2394 3013 2401
rect 3155 2412 3158 2415
rect 3026 2404 3029 2408
rect 3036 2404 3039 2408
rect 3036 2400 3045 2404
rect 3057 2403 3060 2408
rect 3082 2404 3085 2408
rect 3026 2394 3029 2400
rect 3036 2394 3039 2400
rect 3057 2399 3058 2403
rect 3062 2399 3065 2402
rect 3084 2400 3085 2404
rect 3100 2403 3103 2408
rect 3132 2408 3143 2411
rect 3155 2409 3163 2412
rect 3057 2394 3060 2399
rect 3082 2394 3085 2400
rect 3132 2402 3135 2408
rect 3155 2403 3158 2409
rect 3167 2404 3170 2407
rect 3178 2407 3181 2421
rect 3205 2416 3208 2421
rect 3220 2423 3223 2433
rect 3250 2429 3253 2433
rect 3286 2429 3289 2433
rect 3189 2412 3190 2415
rect 3194 2412 3197 2415
rect 3236 2412 3239 2415
rect 3178 2404 3186 2407
rect 3205 2407 3208 2412
rect 3100 2394 3103 2399
rect 3178 2399 3181 2404
rect 3186 2400 3190 2404
rect 3213 2408 3224 2411
rect 3236 2409 3244 2412
rect 3130 2393 3135 2398
rect 3002 2381 3003 2385
rect 3027 2382 3028 2386
rect 3074 2381 3075 2385
rect 2879 2374 2955 2378
rect 2959 2374 3014 2378
rect 3018 2374 3039 2378
rect 3043 2374 3070 2378
rect 3074 2374 3103 2378
rect 3139 2371 3142 2399
rect 3169 2371 3172 2395
rect 3196 2371 3199 2403
rect 3213 2402 3216 2408
rect 3236 2403 3239 2409
rect 3248 2404 3251 2407
rect 3259 2407 3262 2421
rect 3295 2416 3298 2421
rect 3310 2423 3313 2433
rect 3340 2429 3343 2433
rect 3284 2412 3287 2415
rect 3326 2412 3329 2415
rect 3259 2404 3268 2407
rect 3295 2407 3298 2412
rect 3259 2399 3262 2404
rect 3211 2393 3216 2398
rect 3220 2371 3223 2399
rect 3302 2410 3314 2411
rect 3306 2408 3314 2410
rect 3326 2409 3334 2412
rect 3326 2403 3329 2409
rect 3338 2404 3341 2407
rect 3349 2407 3352 2421
rect 3349 2404 3369 2407
rect 3250 2371 3253 2395
rect 3286 2371 3289 2403
rect 3349 2399 3352 2404
rect 3373 2403 4228 2407
rect 3310 2371 3313 2399
rect 3340 2371 3343 2395
rect 1922 2367 1996 2371
rect 2000 2367 2002 2371
rect 2006 2367 2010 2371
rect 2014 2367 2028 2371
rect 2032 2367 2037 2371
rect 2041 2367 2046 2371
rect 2050 2367 2069 2371
rect 2073 2367 2103 2371
rect 2107 2367 2118 2371
rect 2122 2367 2146 2371
rect 2150 2367 2163 2371
rect 2167 2367 2187 2371
rect 2191 2367 2241 2371
rect 2248 2367 2268 2371
rect 2272 2367 2322 2371
rect 2326 2367 2358 2371
rect 2362 2367 2412 2371
rect 2867 2367 2941 2371
rect 2945 2367 2947 2371
rect 2951 2367 2955 2371
rect 2959 2367 2973 2371
rect 2977 2367 2982 2371
rect 2986 2367 2991 2371
rect 2995 2367 3014 2371
rect 3018 2367 3048 2371
rect 3052 2367 3063 2371
rect 3067 2367 3091 2371
rect 3095 2367 3108 2371
rect 3112 2367 3132 2371
rect 3136 2367 3186 2371
rect 3193 2367 3213 2371
rect 3217 2367 3267 2371
rect 3271 2367 3303 2371
rect 3307 2367 3357 2371
rect 1934 2360 2010 2364
rect 2014 2360 2069 2364
rect 2073 2360 2094 2364
rect 2098 2360 2125 2364
rect 2129 2360 2158 2364
rect 2057 2353 2058 2357
rect 2082 2352 2083 2356
rect 2129 2353 2130 2357
rect 2005 2339 2008 2344
rect 2012 2339 2015 2344
rect 1995 2336 1997 2339
rect 2005 2336 2015 2339
rect 2005 2330 2008 2336
rect 2012 2330 2015 2336
rect 2021 2338 2024 2344
rect 2037 2339 2040 2344
rect 2021 2334 2023 2338
rect 2027 2334 2029 2338
rect 2037 2337 2043 2339
rect 2047 2337 2048 2339
rect 2037 2335 2048 2337
rect 2065 2337 2068 2344
rect 2021 2330 2024 2334
rect 2037 2330 2040 2335
rect 2066 2333 2068 2337
rect 2065 2330 2068 2333
rect 2081 2338 2084 2344
rect 2091 2338 2094 2344
rect 2112 2339 2115 2344
rect 2091 2334 2100 2338
rect 2112 2335 2113 2339
rect 2117 2336 2120 2339
rect 2137 2338 2140 2344
rect 2155 2339 2158 2344
rect 2194 2345 2197 2367
rect 2275 2345 2278 2367
rect 2365 2345 2368 2367
rect 2879 2360 2955 2364
rect 2959 2360 3014 2364
rect 3018 2360 3039 2364
rect 3043 2360 3070 2364
rect 3074 2360 3103 2364
rect 3002 2353 3003 2357
rect 3027 2352 3028 2356
rect 3074 2353 3075 2357
rect 2081 2330 2084 2334
rect 2091 2330 2094 2334
rect 2112 2330 2115 2335
rect 2139 2334 2140 2338
rect 2137 2330 2140 2334
rect 2155 2330 2158 2335
rect 2185 2332 2190 2337
rect 2194 2333 2195 2336
rect 2210 2335 2213 2341
rect 2210 2332 2218 2335
rect 2265 2332 2270 2337
rect 2274 2333 2276 2336
rect 2291 2335 2294 2341
rect 2291 2332 2299 2335
rect 2358 2333 2366 2336
rect 2381 2335 2384 2341
rect 2950 2339 2953 2344
rect 2957 2339 2960 2344
rect 2940 2336 2942 2339
rect 2381 2332 2389 2335
rect 2950 2336 2960 2339
rect 2210 2329 2213 2332
rect 2291 2329 2294 2332
rect 2381 2329 2384 2332
rect 2950 2330 2953 2336
rect 2065 2315 2068 2319
rect 2092 2315 2093 2319
rect 2137 2315 2139 2319
rect 2957 2330 2960 2336
rect 2966 2338 2969 2344
rect 2982 2339 2985 2344
rect 2966 2334 2968 2338
rect 2972 2334 2974 2338
rect 2982 2337 2988 2339
rect 2992 2337 2993 2339
rect 2982 2335 2993 2337
rect 3010 2337 3013 2344
rect 2966 2330 2969 2334
rect 2982 2330 2985 2335
rect 3011 2333 3013 2337
rect 3010 2330 3013 2333
rect 3026 2338 3029 2344
rect 3036 2338 3039 2344
rect 3057 2339 3060 2344
rect 3036 2334 3045 2338
rect 3057 2335 3058 2339
rect 3062 2336 3065 2339
rect 3082 2338 3085 2344
rect 3100 2339 3103 2344
rect 3139 2345 3142 2367
rect 3220 2345 3223 2367
rect 3310 2345 3313 2367
rect 4240 2342 4324 2355
rect 3026 2330 3029 2334
rect 3036 2330 3039 2334
rect 3057 2330 3060 2335
rect 3084 2334 3085 2338
rect 3082 2330 3085 2334
rect 3100 2330 3103 2335
rect 3130 2332 3135 2337
rect 3139 2333 3140 2336
rect 3155 2335 3158 2341
rect 3155 2332 3163 2335
rect 3210 2332 3215 2337
rect 3219 2333 3221 2336
rect 3236 2335 3239 2341
rect 3236 2332 3244 2335
rect 3303 2333 3311 2336
rect 3326 2335 3329 2341
rect 3326 2332 3334 2335
rect 3155 2329 3158 2332
rect 3236 2329 3239 2332
rect 3326 2329 3329 2332
rect 1946 2308 2022 2312
rect 2026 2308 2053 2312
rect 2057 2308 2075 2312
rect 2079 2308 2140 2312
rect 2144 2308 2158 2312
rect 2194 2305 2197 2321
rect 2275 2305 2278 2321
rect 2365 2305 2368 2321
rect 3010 2315 3013 2319
rect 3037 2315 3038 2319
rect 3082 2315 3084 2319
rect 2891 2308 2967 2312
rect 2971 2308 2998 2312
rect 3002 2308 3020 2312
rect 3024 2308 3085 2312
rect 3089 2308 3103 2312
rect 3139 2305 3142 2321
rect 3220 2305 3223 2321
rect 3310 2305 3313 2321
rect 1910 2301 1995 2305
rect 1999 2301 2011 2305
rect 2015 2301 2029 2305
rect 2033 2301 2040 2305
rect 2044 2301 2046 2305
rect 2050 2301 2065 2305
rect 2069 2301 2102 2305
rect 2106 2301 2107 2305
rect 2111 2301 2119 2305
rect 2123 2301 2147 2305
rect 2151 2301 2163 2305
rect 2167 2301 2187 2305
rect 2191 2301 2241 2305
rect 2245 2301 2268 2305
rect 2272 2301 2358 2305
rect 2362 2301 2416 2305
rect 2855 2301 2940 2305
rect 2944 2301 2956 2305
rect 2960 2301 2974 2305
rect 2978 2301 2985 2305
rect 2989 2301 2991 2305
rect 2995 2301 3010 2305
rect 3014 2301 3047 2305
rect 3051 2301 3052 2305
rect 3056 2301 3064 2305
rect 3068 2301 3092 2305
rect 3096 2301 3108 2305
rect 3112 2301 3132 2305
rect 3136 2301 3186 2305
rect 3190 2301 3213 2305
rect 3217 2301 3303 2305
rect 3307 2301 3361 2305
rect 1946 2294 2022 2298
rect 2026 2294 2053 2298
rect 2057 2294 2075 2298
rect 2079 2294 2140 2298
rect 2144 2294 2158 2298
rect 2194 2291 2197 2301
rect 2224 2297 2227 2301
rect 2065 2287 2068 2291
rect 2092 2287 2093 2291
rect 2137 2287 2139 2291
rect 1994 2267 1997 2270
rect 2005 2270 2008 2276
rect 2012 2270 2015 2276
rect 2005 2267 2015 2270
rect 2005 2262 2008 2267
rect 2012 2262 2015 2267
rect 2021 2272 2024 2276
rect 2021 2268 2023 2272
rect 2027 2268 2029 2272
rect 2037 2271 2040 2276
rect 2065 2273 2068 2276
rect 2037 2269 2048 2271
rect 2021 2262 2024 2268
rect 2037 2267 2043 2269
rect 2037 2262 2040 2267
rect 2047 2267 2048 2269
rect 2066 2269 2068 2273
rect 2065 2262 2068 2269
rect 2891 2294 2967 2298
rect 2971 2294 2998 2298
rect 3002 2294 3020 2298
rect 3024 2294 3085 2298
rect 3089 2294 3103 2298
rect 3139 2291 3142 2301
rect 3169 2297 3172 2301
rect 2210 2280 2213 2283
rect 2081 2272 2084 2276
rect 2091 2272 2094 2276
rect 2091 2268 2100 2272
rect 2112 2271 2115 2276
rect 2137 2272 2140 2276
rect 2081 2262 2084 2268
rect 2091 2262 2094 2268
rect 2112 2267 2113 2271
rect 2117 2267 2120 2270
rect 2139 2268 2140 2272
rect 2155 2271 2158 2276
rect 2187 2276 2198 2279
rect 2210 2277 2218 2280
rect 2112 2262 2115 2267
rect 2137 2262 2140 2268
rect 2187 2270 2190 2276
rect 2210 2271 2213 2277
rect 2222 2272 2225 2275
rect 2233 2275 2236 2289
rect 3010 2287 3013 2291
rect 3037 2287 3038 2291
rect 3082 2287 3084 2291
rect 2241 2275 2246 2280
rect 2233 2272 2241 2275
rect 2155 2262 2158 2267
rect 2233 2267 2236 2272
rect 2939 2267 2942 2270
rect 2950 2270 2953 2276
rect 2957 2270 2960 2276
rect 2950 2267 2960 2270
rect 2185 2261 2190 2266
rect 1504 2246 1513 2250
rect 1517 2246 1549 2250
rect 1553 2246 1616 2250
rect 1620 2246 1645 2250
rect 1649 2246 1681 2250
rect 1685 2246 1748 2250
rect 1752 2246 1777 2250
rect 1781 2246 1813 2250
rect 1817 2246 1880 2250
rect 1884 2246 1964 2250
rect 2057 2249 2058 2253
rect 2082 2250 2083 2254
rect 2129 2249 2130 2253
rect 1504 2239 1537 2243
rect 1541 2239 1565 2243
rect 1569 2239 1595 2243
rect 1599 2239 1632 2243
rect 1636 2239 1669 2243
rect 1673 2239 1697 2243
rect 1701 2239 1727 2243
rect 1731 2239 1764 2243
rect 1768 2239 1801 2243
rect 1805 2239 1829 2243
rect 1833 2239 1859 2243
rect 1863 2239 1896 2243
rect 1900 2239 1904 2243
rect 1989 2242 2010 2246
rect 2014 2242 2019 2246
rect 2023 2242 2069 2246
rect 2073 2242 2094 2246
rect 2098 2242 2125 2246
rect 2129 2242 2158 2246
rect 2194 2239 2197 2267
rect 2224 2239 2227 2263
rect 2950 2262 2953 2267
rect 2957 2262 2960 2267
rect 2966 2272 2969 2276
rect 2966 2268 2968 2272
rect 2972 2268 2974 2272
rect 2982 2271 2985 2276
rect 3010 2273 3013 2276
rect 2982 2269 2993 2271
rect 2966 2262 2969 2268
rect 2982 2267 2988 2269
rect 2982 2262 2985 2267
rect 2992 2267 2993 2269
rect 3011 2269 3013 2273
rect 3010 2262 3013 2269
rect 3155 2280 3158 2283
rect 3026 2272 3029 2276
rect 3036 2272 3039 2276
rect 3036 2268 3045 2272
rect 3057 2271 3060 2276
rect 3082 2272 3085 2276
rect 3026 2262 3029 2268
rect 3036 2262 3039 2268
rect 3057 2267 3058 2271
rect 3062 2267 3065 2270
rect 3084 2268 3085 2272
rect 3100 2271 3103 2276
rect 3132 2276 3143 2279
rect 3155 2277 3163 2280
rect 3057 2262 3060 2267
rect 3082 2262 3085 2268
rect 3132 2270 3135 2276
rect 3155 2271 3158 2277
rect 3167 2272 3170 2275
rect 3178 2275 3181 2289
rect 3186 2275 3191 2280
rect 3178 2272 3186 2275
rect 3100 2262 3103 2267
rect 3178 2267 3181 2272
rect 3130 2261 3135 2266
rect 2449 2246 2458 2250
rect 2462 2246 2494 2250
rect 2498 2246 2561 2250
rect 2565 2246 2590 2250
rect 2594 2246 2626 2250
rect 2630 2246 2693 2250
rect 2697 2246 2722 2250
rect 2726 2246 2758 2250
rect 2762 2246 2825 2250
rect 2829 2246 2909 2250
rect 3002 2249 3003 2253
rect 3027 2250 3028 2254
rect 3074 2249 3075 2253
rect 2449 2239 2482 2243
rect 2486 2239 2510 2243
rect 2514 2239 2540 2243
rect 2544 2239 2577 2243
rect 2581 2239 2614 2243
rect 2618 2239 2642 2243
rect 2646 2239 2672 2243
rect 2676 2239 2709 2243
rect 2713 2239 2746 2243
rect 2750 2239 2774 2243
rect 2778 2239 2804 2243
rect 2808 2239 2841 2243
rect 2845 2239 2849 2243
rect 2934 2242 2955 2246
rect 2959 2242 2964 2246
rect 2968 2242 3014 2246
rect 3018 2242 3039 2246
rect 3043 2242 3070 2246
rect 3074 2242 3103 2246
rect 3139 2239 3142 2267
rect 3169 2239 3172 2263
rect 1507 2229 1510 2239
rect 1528 2229 1531 2239
rect 1544 2229 1547 2239
rect 1558 2232 1563 2236
rect 1567 2232 1574 2236
rect 1586 2229 1589 2239
rect 1602 2229 1605 2239
rect 1623 2229 1626 2239
rect 1639 2229 1642 2239
rect 1660 2229 1663 2239
rect 1676 2229 1679 2239
rect 1690 2232 1695 2236
rect 1699 2232 1706 2236
rect 1718 2229 1721 2239
rect 1734 2229 1737 2239
rect 1755 2229 1758 2239
rect 1771 2229 1774 2239
rect 1792 2229 1795 2239
rect 1808 2229 1811 2239
rect 1822 2232 1827 2236
rect 1831 2232 1838 2236
rect 1850 2229 1853 2239
rect 1866 2229 1869 2239
rect 1887 2229 1890 2239
rect 1922 2235 1996 2239
rect 2000 2235 2002 2239
rect 2006 2235 2010 2239
rect 2014 2235 2028 2239
rect 2032 2235 2037 2239
rect 2041 2235 2046 2239
rect 2050 2235 2069 2239
rect 2073 2235 2103 2239
rect 2107 2235 2118 2239
rect 2122 2235 2146 2239
rect 2150 2235 2163 2239
rect 2167 2235 2187 2239
rect 2191 2235 2271 2239
rect 2275 2235 2289 2239
rect 2293 2235 2298 2239
rect 2302 2235 2307 2239
rect 2311 2235 2330 2239
rect 2334 2235 2364 2239
rect 2368 2235 2379 2239
rect 2383 2235 2407 2239
rect 2411 2235 2420 2239
rect 1524 2215 1529 2218
rect 1533 2215 1557 2218
rect 1582 2215 1589 2218
rect 1593 2215 1615 2218
rect 1635 2215 1642 2218
rect 1656 2215 1661 2218
rect 1665 2215 1689 2218
rect 1714 2215 1721 2218
rect 1725 2215 1747 2218
rect 1767 2215 1774 2218
rect 1788 2215 1793 2218
rect 1797 2215 1821 2218
rect 1934 2228 2010 2232
rect 2014 2228 2019 2232
rect 2023 2228 2069 2232
rect 2073 2228 2094 2232
rect 2098 2228 2125 2232
rect 2129 2228 2158 2232
rect 1846 2215 1853 2218
rect 1857 2215 1879 2218
rect 2057 2221 2058 2225
rect 2082 2220 2083 2224
rect 2129 2221 2130 2225
rect 1540 2205 1547 2208
rect 1551 2209 1570 2212
rect 1570 2202 1573 2208
rect 1598 2205 1605 2208
rect 1609 2209 1624 2212
rect 1672 2205 1679 2208
rect 1683 2209 1702 2212
rect 1702 2202 1705 2208
rect 1730 2205 1737 2208
rect 1741 2209 1756 2212
rect 1804 2205 1811 2208
rect 1815 2209 1834 2212
rect 1834 2202 1837 2208
rect 1862 2205 1869 2208
rect 1873 2209 1890 2212
rect 2005 2207 2008 2212
rect 2012 2207 2015 2212
rect 1995 2204 1997 2207
rect 2005 2204 2015 2207
rect 2005 2198 2008 2204
rect 1507 2186 1510 2198
rect 1528 2186 1531 2198
rect 1544 2186 1547 2198
rect 1558 2189 1570 2192
rect 1586 2186 1589 2198
rect 1602 2186 1605 2198
rect 1623 2186 1626 2198
rect 1639 2186 1642 2198
rect 1660 2186 1663 2198
rect 1676 2186 1679 2198
rect 1690 2189 1702 2192
rect 1718 2186 1721 2198
rect 1734 2186 1737 2198
rect 1755 2186 1758 2198
rect 1771 2186 1774 2198
rect 1792 2186 1795 2198
rect 1808 2186 1811 2198
rect 1822 2189 1834 2192
rect 1850 2186 1853 2198
rect 1866 2186 1869 2198
rect 1887 2186 1890 2198
rect 2012 2198 2015 2204
rect 2021 2206 2024 2212
rect 2037 2207 2040 2212
rect 2021 2202 2023 2206
rect 2027 2202 2029 2206
rect 2037 2205 2043 2207
rect 2047 2205 2048 2207
rect 2037 2203 2048 2205
rect 2065 2205 2068 2212
rect 2021 2198 2024 2202
rect 2037 2198 2040 2203
rect 2066 2201 2068 2205
rect 2065 2198 2068 2201
rect 2081 2206 2084 2212
rect 2091 2206 2094 2212
rect 2112 2207 2115 2212
rect 2091 2202 2100 2206
rect 2112 2203 2113 2207
rect 2117 2204 2120 2207
rect 2137 2206 2140 2212
rect 2155 2207 2158 2212
rect 2194 2209 2197 2235
rect 2230 2228 2249 2232
rect 2253 2228 2271 2232
rect 2275 2228 2330 2232
rect 2334 2228 2355 2232
rect 2359 2228 2386 2232
rect 2390 2228 2419 2232
rect 2452 2229 2455 2239
rect 2473 2229 2476 2239
rect 2489 2229 2492 2239
rect 2503 2232 2508 2236
rect 2512 2232 2519 2236
rect 2531 2229 2534 2239
rect 2547 2229 2550 2239
rect 2568 2229 2571 2239
rect 2584 2229 2587 2239
rect 2605 2229 2608 2239
rect 2621 2229 2624 2239
rect 2635 2232 2640 2236
rect 2644 2232 2651 2236
rect 2663 2229 2666 2239
rect 2679 2229 2682 2239
rect 2700 2229 2703 2239
rect 2716 2229 2719 2239
rect 2737 2229 2740 2239
rect 2753 2229 2756 2239
rect 2767 2232 2772 2236
rect 2776 2232 2783 2236
rect 2795 2229 2798 2239
rect 2811 2229 2814 2239
rect 2832 2229 2835 2239
rect 2867 2235 2941 2239
rect 2945 2235 2947 2239
rect 2951 2235 2955 2239
rect 2959 2235 2973 2239
rect 2977 2235 2982 2239
rect 2986 2235 2991 2239
rect 2995 2235 3014 2239
rect 3018 2235 3048 2239
rect 3052 2235 3063 2239
rect 3067 2235 3091 2239
rect 3095 2235 3108 2239
rect 3112 2235 3132 2239
rect 3136 2235 3216 2239
rect 3220 2235 3234 2239
rect 3238 2235 3243 2239
rect 3247 2235 3252 2239
rect 3256 2235 3275 2239
rect 3279 2235 3309 2239
rect 3313 2235 3324 2239
rect 3328 2235 3352 2239
rect 3356 2235 3365 2239
rect 2230 2216 2233 2228
rect 2318 2221 2319 2225
rect 2343 2220 2344 2224
rect 2390 2221 2391 2225
rect 2081 2198 2084 2202
rect 2091 2198 2094 2202
rect 2112 2198 2115 2203
rect 2139 2202 2140 2206
rect 2257 2207 2260 2212
rect 2266 2207 2269 2212
rect 2273 2207 2276 2212
rect 2137 2198 2140 2202
rect 2155 2198 2158 2203
rect 2184 2196 2189 2201
rect 2193 2197 2195 2200
rect 2210 2199 2213 2205
rect 2242 2204 2276 2207
rect 2210 2196 2218 2199
rect 2210 2193 2213 2196
rect 1504 2182 1537 2186
rect 1541 2182 1565 2186
rect 1569 2182 1595 2186
rect 1599 2182 1669 2186
rect 1673 2182 1697 2186
rect 1701 2182 1727 2186
rect 1731 2182 1801 2186
rect 1805 2182 1829 2186
rect 1833 2182 1859 2186
rect 1863 2182 1916 2186
rect 2065 2183 2068 2187
rect 2092 2183 2093 2187
rect 2137 2183 2139 2187
rect 2242 2190 2245 2204
rect 2266 2198 2269 2204
rect 2273 2198 2276 2204
rect 2282 2206 2285 2212
rect 2298 2207 2301 2212
rect 2282 2202 2284 2206
rect 2288 2202 2290 2206
rect 2298 2205 2304 2207
rect 2308 2205 2309 2207
rect 2298 2203 2309 2205
rect 2326 2205 2329 2212
rect 2282 2198 2285 2202
rect 2298 2198 2301 2203
rect 2327 2201 2329 2205
rect 2326 2198 2329 2201
rect 2469 2215 2474 2218
rect 2478 2215 2502 2218
rect 2527 2215 2534 2218
rect 2538 2215 2560 2218
rect 2580 2215 2587 2218
rect 2601 2215 2606 2218
rect 2610 2215 2634 2218
rect 2659 2215 2666 2218
rect 2670 2215 2692 2218
rect 2712 2215 2719 2218
rect 2733 2215 2738 2218
rect 2742 2215 2766 2218
rect 2879 2228 2955 2232
rect 2959 2228 2964 2232
rect 2968 2228 3014 2232
rect 3018 2228 3039 2232
rect 3043 2228 3070 2232
rect 3074 2228 3103 2232
rect 2791 2215 2798 2218
rect 2802 2215 2824 2218
rect 3002 2221 3003 2225
rect 3027 2220 3028 2224
rect 3074 2221 3075 2225
rect 2342 2206 2345 2212
rect 2352 2206 2355 2212
rect 2373 2207 2376 2212
rect 2352 2202 2361 2206
rect 2373 2203 2374 2207
rect 2378 2204 2381 2207
rect 2398 2206 2401 2212
rect 2416 2207 2419 2212
rect 2342 2198 2345 2202
rect 2352 2198 2355 2202
rect 2373 2198 2376 2203
rect 2400 2202 2401 2206
rect 2398 2198 2401 2202
rect 2416 2198 2419 2203
rect 2485 2205 2492 2208
rect 2496 2209 2515 2212
rect 2515 2202 2518 2208
rect 2543 2205 2550 2208
rect 2554 2209 2569 2212
rect 2617 2205 2624 2208
rect 2628 2209 2647 2212
rect 2647 2202 2650 2208
rect 2675 2205 2682 2208
rect 2686 2209 2701 2212
rect 2749 2205 2756 2208
rect 2760 2209 2779 2212
rect 2779 2202 2782 2208
rect 2807 2205 2814 2208
rect 2818 2209 2835 2212
rect 2950 2207 2953 2212
rect 2957 2207 2960 2212
rect 2940 2204 2942 2207
rect 2950 2204 2960 2207
rect 2950 2198 2953 2204
rect 1504 2175 1513 2179
rect 1517 2175 1564 2179
rect 1568 2175 1614 2179
rect 1618 2175 1645 2179
rect 1649 2175 1696 2179
rect 1700 2175 1746 2179
rect 1750 2175 1777 2179
rect 1781 2175 1828 2179
rect 1832 2175 1878 2179
rect 1882 2176 1952 2179
rect 2008 2176 2022 2180
rect 2026 2176 2053 2180
rect 2057 2176 2075 2180
rect 2079 2176 2140 2180
rect 2144 2176 2158 2180
rect 2194 2173 2197 2185
rect 2326 2183 2329 2187
rect 2353 2183 2354 2187
rect 2398 2183 2400 2187
rect 2452 2186 2455 2198
rect 2473 2186 2476 2198
rect 2489 2186 2492 2198
rect 2503 2189 2515 2192
rect 2531 2186 2534 2198
rect 2547 2186 2550 2198
rect 2568 2186 2571 2198
rect 2584 2186 2587 2198
rect 2605 2186 2608 2198
rect 2621 2186 2624 2198
rect 2635 2189 2647 2192
rect 2663 2186 2666 2198
rect 2679 2186 2682 2198
rect 2700 2186 2703 2198
rect 2716 2186 2719 2198
rect 2737 2186 2740 2198
rect 2753 2186 2756 2198
rect 2767 2189 2779 2192
rect 2795 2186 2798 2198
rect 2811 2186 2814 2198
rect 2832 2186 2835 2198
rect 2957 2198 2960 2204
rect 2966 2206 2969 2212
rect 2982 2207 2985 2212
rect 2966 2202 2968 2206
rect 2972 2202 2974 2206
rect 2982 2205 2988 2207
rect 2992 2205 2993 2207
rect 2982 2203 2993 2205
rect 3010 2205 3013 2212
rect 2966 2198 2969 2202
rect 2982 2198 2985 2203
rect 3011 2201 3013 2205
rect 3010 2198 3013 2201
rect 3026 2206 3029 2212
rect 3036 2206 3039 2212
rect 3057 2207 3060 2212
rect 3036 2202 3045 2206
rect 3057 2203 3058 2207
rect 3062 2204 3065 2207
rect 3082 2206 3085 2212
rect 3100 2207 3103 2212
rect 3139 2209 3142 2235
rect 3175 2228 3194 2232
rect 3198 2228 3216 2232
rect 3220 2228 3275 2232
rect 3279 2228 3300 2232
rect 3304 2228 3331 2232
rect 3335 2228 3364 2232
rect 3175 2216 3178 2228
rect 3263 2221 3264 2225
rect 3288 2220 3289 2224
rect 3335 2221 3336 2225
rect 3026 2198 3029 2202
rect 3036 2198 3039 2202
rect 3057 2198 3060 2203
rect 3084 2202 3085 2206
rect 3202 2207 3205 2212
rect 3211 2207 3214 2212
rect 3218 2207 3221 2212
rect 3082 2198 3085 2202
rect 3100 2198 3103 2203
rect 3129 2196 3134 2201
rect 3138 2197 3140 2200
rect 3155 2199 3158 2205
rect 3187 2204 3221 2207
rect 3155 2196 3163 2199
rect 3155 2193 3158 2196
rect 2449 2182 2482 2186
rect 2486 2182 2510 2186
rect 2514 2182 2540 2186
rect 2544 2182 2614 2186
rect 2618 2182 2642 2186
rect 2646 2182 2672 2186
rect 2676 2182 2746 2186
rect 2750 2182 2774 2186
rect 2778 2182 2804 2186
rect 2808 2182 2861 2186
rect 3010 2183 3013 2187
rect 3037 2183 3038 2187
rect 3082 2183 3084 2187
rect 3187 2190 3190 2204
rect 3211 2198 3214 2204
rect 3218 2198 3221 2204
rect 3227 2206 3230 2212
rect 3243 2207 3246 2212
rect 3227 2202 3229 2206
rect 3233 2202 3235 2206
rect 3243 2205 3249 2207
rect 3253 2205 3254 2207
rect 3243 2203 3254 2205
rect 3271 2205 3274 2212
rect 3227 2198 3230 2202
rect 3243 2198 3246 2203
rect 3272 2201 3274 2205
rect 3271 2198 3274 2201
rect 3287 2206 3290 2212
rect 3297 2206 3300 2212
rect 3318 2207 3321 2212
rect 3297 2202 3306 2206
rect 3318 2203 3319 2207
rect 3323 2204 3326 2207
rect 3343 2206 3346 2212
rect 3361 2207 3364 2212
rect 3287 2198 3290 2202
rect 3297 2198 3300 2202
rect 3318 2198 3321 2203
rect 3345 2202 3346 2206
rect 3343 2198 3346 2202
rect 3361 2198 3364 2203
rect 2234 2176 2239 2180
rect 2243 2176 2283 2180
rect 2287 2176 2314 2180
rect 2318 2176 2336 2180
rect 2340 2176 2401 2180
rect 2405 2176 2419 2180
rect 2449 2175 2458 2179
rect 2462 2175 2509 2179
rect 2513 2175 2559 2179
rect 2563 2175 2590 2179
rect 2594 2175 2641 2179
rect 2645 2175 2691 2179
rect 2695 2175 2722 2179
rect 2726 2175 2773 2179
rect 2777 2175 2823 2179
rect 2827 2176 2897 2179
rect 2953 2176 2967 2180
rect 2971 2176 2998 2180
rect 3002 2176 3020 2180
rect 3024 2176 3085 2180
rect 3089 2176 3103 2180
rect 3139 2173 3142 2185
rect 3271 2183 3274 2187
rect 3298 2183 3299 2187
rect 3343 2183 3345 2187
rect 3179 2176 3184 2180
rect 3188 2176 3228 2180
rect 3232 2176 3259 2180
rect 3263 2176 3281 2180
rect 3285 2176 3346 2180
rect 3350 2176 3364 2180
rect 1511 2169 1895 2172
rect 1910 2169 1995 2173
rect 1999 2169 2011 2173
rect 2015 2169 2029 2173
rect 2033 2169 2040 2173
rect 2044 2169 2046 2173
rect 2050 2169 2065 2173
rect 2069 2169 2102 2173
rect 2106 2169 2107 2173
rect 2111 2169 2119 2173
rect 2123 2169 2147 2173
rect 2151 2169 2187 2173
rect 2191 2169 2230 2173
rect 2234 2169 2241 2173
rect 2245 2169 2256 2173
rect 2260 2169 2272 2173
rect 2276 2169 2290 2173
rect 2294 2169 2301 2173
rect 2305 2169 2307 2173
rect 2311 2169 2326 2173
rect 2330 2169 2363 2173
rect 2367 2169 2368 2173
rect 2372 2169 2380 2173
rect 2384 2169 2408 2173
rect 2412 2169 2420 2173
rect 2456 2169 2840 2172
rect 2855 2169 2940 2173
rect 2944 2169 2956 2173
rect 2960 2169 2974 2173
rect 2978 2169 2985 2173
rect 2989 2169 2991 2173
rect 2995 2169 3010 2173
rect 3014 2169 3047 2173
rect 3051 2169 3052 2173
rect 3056 2169 3064 2173
rect 3068 2169 3092 2173
rect 3096 2169 3132 2173
rect 3136 2169 3175 2173
rect 3179 2169 3186 2173
rect 3190 2169 3201 2173
rect 3205 2169 3217 2173
rect 3221 2169 3235 2173
rect 3239 2169 3246 2173
rect 3250 2169 3252 2173
rect 3256 2169 3271 2173
rect 3275 2169 3308 2173
rect 3312 2169 3313 2173
rect 3317 2169 3325 2173
rect 3329 2169 3353 2173
rect 3357 2169 3365 2173
rect 1654 2162 1763 2165
rect 1946 2162 2004 2166
rect 2008 2162 2238 2165
rect 2428 2163 2436 2167
rect 2599 2162 2708 2165
rect 2891 2162 2949 2166
rect 2953 2162 3183 2165
rect 3373 2163 3381 2167
rect 1634 2154 1638 2158
rect 1642 2154 1646 2158
rect 1934 2155 2248 2158
rect 1982 2148 2255 2152
rect 2424 2145 2428 2151
rect 2579 2154 2583 2158
rect 2587 2154 2591 2158
rect 2879 2155 3193 2158
rect 2927 2148 3198 2152
rect 3369 2145 3373 2151
rect 1490 2141 1622 2145
rect 1626 2141 1642 2145
rect 1658 2141 2567 2145
rect 2571 2141 2587 2145
rect 2603 2141 3461 2145
rect 1650 2134 1895 2137
rect 1970 2134 2296 2138
rect 2300 2134 2332 2138
rect 2336 2134 2399 2138
rect 2403 2134 2419 2138
rect 2595 2134 2840 2137
rect 2915 2134 3241 2138
rect 3245 2134 3277 2138
rect 3281 2134 3344 2138
rect 3348 2134 3364 2138
rect 1665 2127 1895 2130
rect 1910 2127 2282 2131
rect 2286 2127 2320 2131
rect 2324 2127 2348 2131
rect 2352 2127 2378 2131
rect 2382 2127 2415 2131
rect 1634 2118 1638 2122
rect 1642 2118 1646 2122
rect 2290 2117 2293 2127
rect 2311 2117 2314 2127
rect 2327 2117 2330 2127
rect 2341 2120 2346 2124
rect 2350 2120 2357 2124
rect 2369 2117 2372 2127
rect 2385 2117 2388 2127
rect 2406 2117 2409 2127
rect 2610 2127 2840 2130
rect 2855 2127 3227 2131
rect 3231 2127 3265 2131
rect 3269 2127 3293 2131
rect 3297 2127 3323 2131
rect 3327 2127 3360 2131
rect 2579 2118 2583 2122
rect 2587 2118 2591 2122
rect 3235 2117 3238 2127
rect 3256 2117 3259 2127
rect 3272 2117 3275 2127
rect 3286 2120 3291 2124
rect 3295 2120 3302 2124
rect 3314 2117 3317 2127
rect 3330 2117 3333 2127
rect 3351 2117 3354 2127
rect 1654 2111 1764 2114
rect 1504 2104 1513 2108
rect 1517 2104 1549 2108
rect 1553 2104 1616 2108
rect 1620 2104 1645 2108
rect 1649 2104 1681 2108
rect 1685 2104 1748 2108
rect 1752 2104 1777 2108
rect 1781 2104 1813 2108
rect 1817 2104 1880 2108
rect 1884 2104 1964 2108
rect 1504 2097 1537 2101
rect 1541 2097 1565 2101
rect 1569 2097 1595 2101
rect 1599 2097 1632 2101
rect 1636 2097 1669 2101
rect 1673 2097 1697 2101
rect 1701 2097 1727 2101
rect 1731 2097 1764 2101
rect 1768 2097 1801 2101
rect 1805 2097 1829 2101
rect 1833 2097 1859 2101
rect 1863 2097 1896 2101
rect 1900 2097 1904 2101
rect 2307 2103 2312 2106
rect 2316 2103 2340 2106
rect 2599 2111 2709 2114
rect 2365 2103 2372 2106
rect 2376 2103 2398 2106
rect 2449 2104 2458 2108
rect 2462 2104 2494 2108
rect 2498 2104 2561 2108
rect 2565 2104 2590 2108
rect 2594 2104 2626 2108
rect 2630 2104 2693 2108
rect 2697 2104 2722 2108
rect 2726 2104 2758 2108
rect 2762 2104 2825 2108
rect 2829 2104 2909 2108
rect 1507 2087 1510 2097
rect 1528 2087 1531 2097
rect 1544 2087 1547 2097
rect 1558 2090 1563 2094
rect 1567 2090 1574 2094
rect 1586 2087 1589 2097
rect 1602 2087 1605 2097
rect 1623 2087 1626 2097
rect 1639 2087 1642 2097
rect 1660 2087 1663 2097
rect 1676 2087 1679 2097
rect 1690 2090 1695 2094
rect 1699 2090 1706 2094
rect 1718 2087 1721 2097
rect 1734 2087 1737 2097
rect 1755 2087 1758 2097
rect 1771 2087 1774 2097
rect 1792 2087 1795 2097
rect 1808 2087 1811 2097
rect 1822 2090 1827 2094
rect 1831 2090 1838 2094
rect 1850 2087 1853 2097
rect 1866 2087 1869 2097
rect 1887 2087 1890 2097
rect 2323 2093 2330 2096
rect 2334 2097 2353 2100
rect 1524 2073 1529 2076
rect 1533 2073 1557 2076
rect 1582 2073 1589 2076
rect 1593 2073 1615 2076
rect 1635 2073 1642 2076
rect 1656 2073 1661 2076
rect 1665 2073 1689 2076
rect 1714 2073 1721 2076
rect 1725 2073 1747 2076
rect 1767 2073 1774 2076
rect 1788 2073 1793 2076
rect 1797 2073 1821 2076
rect 1846 2073 1853 2076
rect 1857 2073 1879 2076
rect 2353 2090 2356 2096
rect 2381 2093 2388 2096
rect 2392 2097 2407 2100
rect 2449 2097 2482 2101
rect 2486 2097 2510 2101
rect 2514 2097 2540 2101
rect 2544 2097 2577 2101
rect 2581 2097 2614 2101
rect 2618 2097 2642 2101
rect 2646 2097 2672 2101
rect 2676 2097 2709 2101
rect 2713 2097 2746 2101
rect 2750 2097 2774 2101
rect 2778 2097 2804 2101
rect 2808 2097 2841 2101
rect 2845 2097 2849 2101
rect 3252 2103 3257 2106
rect 3261 2103 3285 2106
rect 3310 2103 3317 2106
rect 3321 2103 3343 2106
rect 2452 2087 2455 2097
rect 2473 2087 2476 2097
rect 2489 2087 2492 2097
rect 2503 2090 2508 2094
rect 2512 2090 2519 2094
rect 2531 2087 2534 2097
rect 2547 2087 2550 2097
rect 2568 2087 2571 2097
rect 2584 2087 2587 2097
rect 2605 2087 2608 2097
rect 2621 2087 2624 2097
rect 2635 2090 2640 2094
rect 2644 2090 2651 2094
rect 2663 2087 2666 2097
rect 2679 2087 2682 2097
rect 2700 2087 2703 2097
rect 2716 2087 2719 2097
rect 2737 2087 2740 2097
rect 2753 2087 2756 2097
rect 2767 2090 2772 2094
rect 2776 2090 2783 2094
rect 2795 2087 2798 2097
rect 2811 2087 2814 2097
rect 2832 2087 2835 2097
rect 3268 2093 3275 2096
rect 3279 2097 3298 2100
rect 2290 2074 2293 2086
rect 2311 2074 2314 2086
rect 2327 2074 2330 2086
rect 2341 2077 2353 2080
rect 2369 2074 2372 2086
rect 2385 2074 2388 2086
rect 2406 2074 2409 2086
rect 1540 2063 1547 2066
rect 1551 2067 1570 2070
rect 1570 2060 1573 2066
rect 1598 2063 1605 2066
rect 1609 2067 1624 2070
rect 1672 2063 1679 2066
rect 1683 2067 1702 2070
rect 1702 2060 1705 2066
rect 1730 2063 1737 2066
rect 1741 2067 1756 2070
rect 1804 2063 1811 2066
rect 1815 2067 1834 2070
rect 1834 2060 1837 2066
rect 1862 2063 1869 2066
rect 1873 2067 1890 2070
rect 1922 2070 2320 2074
rect 2324 2070 2348 2074
rect 2352 2070 2378 2074
rect 2382 2070 2419 2074
rect 2469 2073 2474 2076
rect 2478 2073 2502 2076
rect 2527 2073 2534 2076
rect 2538 2073 2560 2076
rect 2580 2073 2587 2076
rect 2601 2073 2606 2076
rect 2610 2073 2634 2076
rect 2659 2073 2666 2076
rect 2670 2073 2692 2076
rect 2712 2073 2719 2076
rect 2733 2073 2738 2076
rect 2742 2073 2766 2076
rect 2791 2073 2798 2076
rect 2802 2073 2824 2076
rect 3298 2090 3301 2096
rect 3326 2093 3333 2096
rect 3337 2097 3352 2100
rect 3235 2074 3238 2086
rect 3256 2074 3259 2086
rect 3272 2074 3275 2086
rect 3286 2077 3298 2080
rect 3314 2074 3317 2086
rect 3330 2074 3333 2086
rect 3351 2074 3354 2086
rect 1958 2063 2296 2067
rect 2300 2063 2347 2067
rect 2351 2063 2397 2067
rect 2401 2063 2419 2067
rect 2485 2063 2492 2066
rect 2496 2067 2515 2070
rect 1507 2044 1510 2056
rect 1528 2044 1531 2056
rect 1544 2044 1547 2056
rect 1558 2047 1570 2050
rect 1586 2044 1589 2056
rect 1602 2044 1605 2056
rect 1623 2044 1626 2056
rect 1639 2044 1642 2056
rect 1660 2044 1663 2056
rect 1676 2044 1679 2056
rect 1690 2047 1702 2050
rect 1718 2044 1721 2056
rect 1734 2044 1737 2056
rect 1755 2044 1758 2056
rect 1771 2044 1774 2056
rect 1792 2044 1795 2056
rect 1808 2044 1811 2056
rect 1822 2047 1834 2050
rect 1850 2044 1853 2056
rect 1866 2044 1869 2056
rect 1887 2044 1890 2056
rect 2293 2056 2414 2059
rect 2515 2060 2518 2066
rect 2543 2063 2550 2066
rect 2554 2067 2569 2070
rect 2617 2063 2624 2066
rect 2628 2067 2647 2070
rect 2647 2060 2650 2066
rect 2675 2063 2682 2066
rect 2686 2067 2701 2070
rect 2749 2063 2756 2066
rect 2760 2067 2779 2070
rect 2779 2060 2782 2066
rect 2807 2063 2814 2066
rect 2818 2067 2835 2070
rect 2867 2070 3265 2074
rect 3269 2070 3293 2074
rect 3297 2070 3323 2074
rect 3327 2070 3364 2074
rect 2903 2063 3241 2067
rect 3245 2063 3292 2067
rect 3296 2063 3342 2067
rect 3346 2063 3364 2067
rect 1970 2048 2296 2052
rect 2300 2048 2332 2052
rect 2336 2048 2399 2052
rect 2403 2048 2419 2052
rect 1504 2040 1537 2044
rect 1541 2040 1565 2044
rect 1569 2040 1595 2044
rect 1599 2040 1669 2044
rect 1673 2040 1697 2044
rect 1701 2040 1727 2044
rect 1731 2040 1801 2044
rect 1805 2040 1829 2044
rect 1833 2040 1859 2044
rect 1863 2040 1916 2044
rect 2286 2041 2320 2045
rect 2324 2041 2348 2045
rect 2352 2041 2378 2045
rect 2382 2041 2415 2045
rect 2452 2044 2455 2056
rect 2473 2044 2476 2056
rect 2489 2044 2492 2056
rect 2503 2047 2515 2050
rect 2531 2044 2534 2056
rect 2547 2044 2550 2056
rect 2568 2044 2571 2056
rect 2584 2044 2587 2056
rect 2605 2044 2608 2056
rect 2621 2044 2624 2056
rect 2635 2047 2647 2050
rect 2663 2044 2666 2056
rect 2679 2044 2682 2056
rect 2700 2044 2703 2056
rect 2716 2044 2719 2056
rect 2737 2044 2740 2056
rect 2753 2044 2756 2056
rect 2767 2047 2779 2050
rect 2795 2044 2798 2056
rect 2811 2044 2814 2056
rect 2832 2044 2835 2056
rect 3238 2056 3359 2059
rect 2915 2048 3241 2052
rect 3245 2048 3277 2052
rect 3281 2048 3344 2052
rect 3348 2048 3364 2052
rect 1504 2033 1513 2037
rect 1517 2033 1564 2037
rect 1568 2033 1614 2037
rect 1618 2033 1645 2037
rect 1649 2033 1696 2037
rect 1700 2033 1746 2037
rect 1750 2033 1777 2037
rect 1781 2033 1828 2037
rect 1832 2033 1878 2037
rect 1882 2033 1952 2037
rect 2290 2031 2293 2041
rect 2311 2031 2314 2041
rect 2327 2031 2330 2041
rect 2341 2034 2346 2038
rect 2350 2034 2357 2038
rect 2369 2031 2372 2041
rect 2385 2031 2388 2041
rect 2406 2031 2409 2041
rect 2449 2040 2482 2044
rect 2486 2040 2510 2044
rect 2514 2040 2540 2044
rect 2544 2040 2614 2044
rect 2618 2040 2642 2044
rect 2646 2040 2672 2044
rect 2676 2040 2746 2044
rect 2750 2040 2774 2044
rect 2778 2040 2804 2044
rect 2808 2040 2861 2044
rect 3231 2041 3265 2045
rect 3269 2041 3293 2045
rect 3297 2041 3323 2045
rect 3327 2041 3360 2045
rect 2449 2033 2458 2037
rect 2462 2033 2509 2037
rect 2513 2033 2559 2037
rect 2563 2033 2590 2037
rect 2594 2033 2641 2037
rect 2645 2033 2691 2037
rect 2695 2033 2722 2037
rect 2726 2033 2773 2037
rect 2777 2033 2823 2037
rect 2827 2033 2897 2037
rect 3235 2031 3238 2041
rect 3256 2031 3259 2041
rect 3272 2031 3275 2041
rect 3286 2034 3291 2038
rect 3295 2034 3302 2038
rect 3314 2031 3317 2041
rect 3330 2031 3333 2041
rect 3351 2031 3354 2041
rect 1510 2026 1895 2029
rect 1504 2018 1513 2022
rect 1517 2018 1549 2022
rect 1553 2018 1616 2022
rect 1620 2018 1645 2022
rect 1649 2018 1681 2022
rect 1685 2018 1748 2022
rect 1752 2018 1777 2022
rect 1781 2018 1813 2022
rect 1817 2018 1880 2022
rect 1884 2018 1964 2022
rect 1504 2011 1537 2015
rect 1541 2011 1565 2015
rect 1569 2011 1595 2015
rect 1599 2011 1632 2015
rect 1636 2011 1669 2015
rect 1673 2011 1697 2015
rect 1701 2011 1727 2015
rect 1731 2011 1764 2015
rect 1768 2011 1801 2015
rect 1805 2011 1829 2015
rect 1833 2011 1859 2015
rect 1863 2011 1896 2015
rect 1900 2011 1904 2015
rect 2307 2017 2312 2020
rect 2316 2017 2340 2020
rect 2455 2026 2840 2029
rect 2365 2017 2372 2020
rect 2376 2017 2398 2020
rect 2449 2018 2458 2022
rect 2462 2018 2494 2022
rect 2498 2018 2561 2022
rect 2565 2018 2590 2022
rect 2594 2018 2626 2022
rect 2630 2018 2693 2022
rect 2697 2018 2722 2022
rect 2726 2018 2758 2022
rect 2762 2018 2825 2022
rect 2829 2018 2909 2022
rect 1507 2001 1510 2011
rect 1528 2001 1531 2011
rect 1544 2001 1547 2011
rect 1558 2004 1563 2008
rect 1567 2004 1574 2008
rect 1586 2001 1589 2011
rect 1602 2001 1605 2011
rect 1623 2001 1626 2011
rect 1639 2001 1642 2011
rect 1660 2001 1663 2011
rect 1676 2001 1679 2011
rect 1690 2004 1695 2008
rect 1699 2004 1706 2008
rect 1718 2001 1721 2011
rect 1734 2001 1737 2011
rect 1755 2001 1758 2011
rect 1771 2001 1774 2011
rect 1792 2001 1795 2011
rect 1808 2001 1811 2011
rect 1822 2004 1827 2008
rect 1831 2004 1838 2008
rect 1850 2001 1853 2011
rect 1866 2001 1869 2011
rect 1887 2001 1890 2011
rect 2323 2007 2330 2010
rect 2334 2011 2353 2014
rect 1524 1987 1529 1990
rect 1533 1987 1557 1990
rect 1582 1987 1589 1990
rect 1593 1987 1615 1990
rect 1635 1987 1642 1990
rect 1656 1987 1661 1990
rect 1665 1987 1689 1990
rect 1714 1987 1721 1990
rect 1725 1987 1747 1990
rect 1767 1987 1774 1990
rect 1788 1987 1793 1990
rect 1797 1987 1821 1990
rect 1846 1987 1853 1990
rect 1857 1987 1879 1990
rect 2353 2004 2356 2010
rect 2381 2007 2388 2010
rect 2392 2011 2407 2014
rect 2418 2009 2429 2013
rect 2449 2011 2482 2015
rect 2486 2011 2510 2015
rect 2514 2011 2540 2015
rect 2544 2011 2577 2015
rect 2581 2011 2614 2015
rect 2618 2011 2642 2015
rect 2646 2011 2672 2015
rect 2676 2011 2709 2015
rect 2713 2011 2746 2015
rect 2750 2011 2774 2015
rect 2778 2011 2804 2015
rect 2808 2011 2841 2015
rect 2845 2011 2849 2015
rect 3252 2017 3257 2020
rect 3261 2017 3285 2020
rect 3310 2017 3317 2020
rect 3321 2017 3343 2020
rect 2452 2001 2455 2011
rect 2473 2001 2476 2011
rect 2489 2001 2492 2011
rect 2503 2004 2508 2008
rect 2512 2004 2519 2008
rect 2531 2001 2534 2011
rect 2547 2001 2550 2011
rect 2568 2001 2571 2011
rect 2584 2001 2587 2011
rect 2605 2001 2608 2011
rect 2621 2001 2624 2011
rect 2635 2004 2640 2008
rect 2644 2004 2651 2008
rect 2663 2001 2666 2011
rect 2679 2001 2682 2011
rect 2700 2001 2703 2011
rect 2716 2001 2719 2011
rect 2737 2001 2740 2011
rect 2753 2001 2756 2011
rect 2767 2004 2772 2008
rect 2776 2004 2783 2008
rect 2795 2001 2798 2011
rect 2811 2001 2814 2011
rect 2832 2001 2835 2011
rect 3268 2007 3275 2010
rect 3279 2011 3298 2014
rect 2290 1988 2293 2000
rect 2311 1988 2314 2000
rect 2327 1988 2330 2000
rect 2341 1991 2353 1994
rect 2369 1988 2372 2000
rect 2385 1988 2388 2000
rect 2406 1988 2409 2000
rect 1540 1977 1547 1980
rect 1551 1981 1570 1984
rect 1570 1974 1573 1980
rect 1598 1977 1605 1980
rect 1609 1981 1624 1984
rect 1672 1977 1679 1980
rect 1683 1981 1702 1984
rect 1702 1974 1705 1980
rect 1730 1977 1737 1980
rect 1741 1981 1756 1984
rect 1804 1977 1811 1980
rect 1815 1981 1834 1984
rect 1834 1974 1837 1980
rect 1862 1977 1869 1980
rect 1873 1981 1890 1984
rect 1922 1984 2320 1988
rect 2324 1984 2348 1988
rect 2352 1984 2378 1988
rect 2382 1984 2419 1988
rect 2469 1987 2474 1990
rect 2478 1987 2502 1990
rect 2527 1987 2534 1990
rect 2538 1987 2560 1990
rect 2580 1987 2587 1990
rect 2601 1987 2606 1990
rect 2610 1987 2634 1990
rect 2659 1987 2666 1990
rect 2670 1987 2692 1990
rect 2712 1987 2719 1990
rect 2733 1987 2738 1990
rect 2742 1987 2766 1990
rect 2791 1987 2798 1990
rect 2802 1987 2824 1990
rect 3298 2004 3301 2010
rect 3326 2007 3333 2010
rect 3337 2011 3352 2014
rect 3363 2009 3374 2013
rect 3235 1988 3238 2000
rect 3256 1988 3259 2000
rect 3272 1988 3275 2000
rect 3286 1991 3298 1994
rect 3314 1988 3317 2000
rect 3330 1988 3333 2000
rect 3351 1988 3354 2000
rect 1958 1977 2296 1981
rect 2300 1977 2347 1981
rect 2351 1977 2397 1981
rect 2401 1977 2419 1981
rect 2485 1977 2492 1980
rect 2496 1981 2515 1984
rect 2515 1974 2518 1980
rect 2543 1977 2550 1980
rect 2554 1981 2569 1984
rect 2617 1977 2624 1980
rect 2628 1981 2647 1984
rect 2647 1974 2650 1980
rect 2675 1977 2682 1980
rect 2686 1981 2701 1984
rect 2749 1977 2756 1980
rect 2760 1981 2779 1984
rect 2779 1974 2782 1980
rect 2807 1977 2814 1980
rect 2818 1981 2835 1984
rect 2867 1984 3265 1988
rect 3269 1984 3293 1988
rect 3297 1984 3323 1988
rect 3327 1984 3364 1988
rect 2903 1977 3241 1981
rect 3245 1977 3292 1981
rect 3296 1977 3342 1981
rect 3346 1977 3364 1981
rect 1507 1958 1510 1970
rect 1528 1958 1531 1970
rect 1544 1958 1547 1970
rect 1558 1961 1570 1964
rect 1586 1958 1589 1970
rect 1602 1958 1605 1970
rect 1623 1958 1626 1970
rect 1639 1958 1642 1970
rect 1660 1958 1663 1970
rect 1676 1958 1679 1970
rect 1690 1961 1702 1964
rect 1718 1958 1721 1970
rect 1734 1958 1737 1970
rect 1755 1958 1758 1970
rect 1771 1958 1774 1970
rect 1792 1958 1795 1970
rect 1808 1958 1811 1970
rect 1822 1961 1834 1964
rect 1850 1958 1853 1970
rect 1866 1958 1869 1970
rect 1887 1958 1890 1970
rect 2452 1958 2455 1970
rect 2473 1958 2476 1970
rect 2489 1958 2492 1970
rect 2503 1961 2515 1964
rect 2531 1958 2534 1970
rect 2547 1958 2550 1970
rect 2568 1958 2571 1970
rect 2584 1958 2587 1970
rect 2605 1958 2608 1970
rect 2621 1958 2624 1970
rect 2635 1961 2647 1964
rect 2663 1958 2666 1970
rect 2679 1958 2682 1970
rect 2700 1958 2703 1970
rect 2716 1958 2719 1970
rect 2737 1958 2740 1970
rect 2753 1958 2756 1970
rect 2767 1961 2779 1964
rect 2795 1958 2798 1970
rect 2811 1958 2814 1970
rect 2832 1958 2835 1970
rect 1504 1954 1537 1958
rect 1541 1954 1565 1958
rect 1569 1954 1595 1958
rect 1599 1954 1669 1958
rect 1673 1954 1697 1958
rect 1701 1954 1727 1958
rect 1731 1954 1801 1958
rect 1805 1954 1829 1958
rect 1833 1954 1859 1958
rect 1863 1954 1916 1958
rect 2449 1954 2482 1958
rect 2486 1954 2510 1958
rect 2514 1954 2540 1958
rect 2544 1954 2614 1958
rect 2618 1954 2642 1958
rect 2646 1954 2672 1958
rect 2676 1954 2746 1958
rect 2750 1954 2774 1958
rect 2778 1954 2804 1958
rect 2808 1954 2861 1958
rect 1504 1947 1513 1951
rect 1517 1947 1564 1951
rect 1568 1947 1614 1951
rect 1618 1947 1645 1951
rect 1649 1947 1696 1951
rect 1700 1947 1746 1951
rect 1750 1947 1777 1951
rect 1781 1947 1828 1951
rect 1832 1947 1878 1951
rect 1882 1947 1952 1951
rect 2449 1947 2458 1951
rect 2462 1947 2509 1951
rect 2513 1947 2559 1951
rect 2563 1947 2590 1951
rect 2594 1947 2641 1951
rect 2645 1947 2691 1951
rect 2695 1947 2722 1951
rect 2726 1947 2773 1951
rect 2777 1947 2823 1951
rect 2827 1947 2897 1951
rect 1510 1941 1895 1944
rect 2455 1941 2840 1944
rect 1635 1934 1739 1937
rect 2580 1934 2684 1937
rect 1751 1926 1755 1930
rect 1759 1926 1763 1930
rect 2696 1926 2700 1930
rect 2704 1926 2708 1930
rect 1487 1915 1739 1919
rect 1743 1915 1759 1919
rect 1775 1915 2436 1919
rect 2440 1915 2684 1919
rect 2688 1915 2704 1919
rect 2720 1915 3381 1919
rect 3385 1915 3468 1919
rect 1767 1908 1895 1911
rect 2712 1908 2840 1911
rect 1782 1901 1895 1904
rect 2727 1901 2840 1904
rect 1751 1892 1755 1896
rect 1759 1892 1763 1896
rect 2696 1892 2700 1896
rect 2704 1892 2708 1896
rect 1635 1885 1739 1888
rect 2580 1885 2684 1888
rect 1504 1878 1513 1882
rect 1517 1878 1549 1882
rect 1553 1878 1616 1882
rect 1620 1878 1645 1882
rect 1649 1878 1681 1882
rect 1685 1878 1748 1882
rect 1752 1878 1777 1882
rect 1781 1878 1813 1882
rect 1817 1878 1880 1882
rect 1884 1878 1964 1882
rect 2449 1878 2458 1882
rect 2462 1878 2494 1882
rect 2498 1878 2561 1882
rect 2565 1878 2590 1882
rect 2594 1878 2626 1882
rect 2630 1878 2693 1882
rect 2697 1878 2722 1882
rect 2726 1878 2758 1882
rect 2762 1878 2825 1882
rect 2829 1878 2909 1882
rect 1504 1871 1537 1875
rect 1541 1871 1565 1875
rect 1569 1871 1595 1875
rect 1599 1871 1632 1875
rect 1636 1871 1669 1875
rect 1673 1871 1697 1875
rect 1701 1871 1727 1875
rect 1731 1871 1764 1875
rect 1768 1871 1801 1875
rect 1805 1871 1829 1875
rect 1833 1871 1859 1875
rect 1863 1871 1896 1875
rect 1900 1871 1904 1875
rect 2449 1871 2482 1875
rect 2486 1871 2510 1875
rect 2514 1871 2540 1875
rect 2544 1871 2577 1875
rect 2581 1871 2614 1875
rect 2618 1871 2642 1875
rect 2646 1871 2672 1875
rect 2676 1871 2709 1875
rect 2713 1871 2746 1875
rect 2750 1871 2774 1875
rect 2778 1871 2804 1875
rect 2808 1871 2841 1875
rect 2845 1871 2849 1875
rect 1507 1861 1510 1871
rect 1528 1861 1531 1871
rect 1544 1861 1547 1871
rect 1558 1864 1563 1868
rect 1567 1864 1574 1868
rect 1586 1861 1589 1871
rect 1602 1861 1605 1871
rect 1623 1861 1626 1871
rect 1639 1861 1642 1871
rect 1660 1861 1663 1871
rect 1676 1861 1679 1871
rect 1690 1864 1695 1868
rect 1699 1864 1706 1868
rect 1718 1861 1721 1871
rect 1734 1861 1737 1871
rect 1755 1861 1758 1871
rect 1771 1861 1774 1871
rect 1792 1861 1795 1871
rect 1808 1861 1811 1871
rect 1822 1864 1827 1868
rect 1831 1864 1838 1868
rect 1850 1861 1853 1871
rect 1866 1861 1869 1871
rect 1887 1861 1890 1871
rect 2452 1861 2455 1871
rect 2473 1861 2476 1871
rect 2489 1861 2492 1871
rect 2503 1864 2508 1868
rect 2512 1864 2519 1868
rect 2531 1861 2534 1871
rect 2547 1861 2550 1871
rect 2568 1861 2571 1871
rect 2584 1861 2587 1871
rect 2605 1861 2608 1871
rect 2621 1861 2624 1871
rect 2635 1864 2640 1868
rect 2644 1864 2651 1868
rect 2663 1861 2666 1871
rect 2679 1861 2682 1871
rect 2700 1861 2703 1871
rect 2716 1861 2719 1871
rect 2737 1861 2740 1871
rect 2753 1861 2756 1871
rect 2767 1864 2772 1868
rect 2776 1864 2783 1868
rect 2795 1861 2798 1871
rect 2811 1861 2814 1871
rect 2832 1861 2835 1871
rect 1524 1847 1529 1850
rect 1533 1847 1557 1850
rect 1582 1847 1589 1850
rect 1593 1847 1615 1850
rect 1635 1847 1642 1850
rect 1656 1847 1661 1850
rect 1665 1847 1689 1850
rect 1714 1847 1721 1850
rect 1725 1847 1747 1850
rect 1767 1847 1774 1850
rect 1788 1847 1793 1850
rect 1797 1847 1821 1850
rect 1846 1847 1853 1850
rect 1857 1847 1879 1850
rect 1540 1837 1547 1840
rect 1551 1841 1570 1844
rect 1570 1834 1573 1840
rect 1598 1837 1605 1840
rect 1609 1841 1624 1844
rect 1672 1837 1679 1840
rect 1683 1841 1702 1844
rect 1702 1834 1705 1840
rect 1730 1837 1737 1840
rect 1741 1841 1756 1844
rect 1804 1837 1811 1840
rect 1815 1841 1834 1844
rect 1834 1834 1837 1840
rect 1862 1837 1869 1840
rect 1873 1841 1890 1844
rect 2469 1847 2474 1850
rect 2478 1847 2502 1850
rect 2527 1847 2534 1850
rect 2538 1847 2560 1850
rect 2580 1847 2587 1850
rect 2601 1847 2606 1850
rect 2610 1847 2634 1850
rect 2659 1847 2666 1850
rect 2670 1847 2692 1850
rect 2712 1847 2719 1850
rect 2733 1847 2738 1850
rect 2742 1847 2766 1850
rect 2791 1847 2798 1850
rect 2802 1847 2824 1850
rect 2485 1837 2492 1840
rect 2496 1841 2515 1844
rect 2515 1834 2518 1840
rect 2543 1837 2550 1840
rect 2554 1841 2569 1844
rect 2617 1837 2624 1840
rect 2628 1841 2647 1844
rect 2647 1834 2650 1840
rect 2675 1837 2682 1840
rect 2686 1841 2701 1844
rect 2749 1837 2756 1840
rect 2760 1841 2779 1844
rect 2779 1834 2782 1840
rect 2807 1837 2814 1840
rect 2818 1841 2835 1844
rect 1507 1818 1510 1830
rect 1528 1818 1531 1830
rect 1544 1818 1547 1830
rect 1558 1821 1570 1824
rect 1586 1818 1589 1830
rect 1602 1818 1605 1830
rect 1623 1818 1626 1830
rect 1639 1818 1642 1830
rect 1660 1818 1663 1830
rect 1676 1818 1679 1830
rect 1690 1821 1702 1824
rect 1718 1818 1721 1830
rect 1734 1818 1737 1830
rect 1755 1818 1758 1830
rect 1771 1818 1774 1830
rect 1792 1818 1795 1830
rect 1808 1818 1811 1830
rect 1822 1821 1834 1824
rect 1850 1818 1853 1830
rect 1866 1818 1869 1830
rect 1887 1818 1890 1830
rect 2452 1818 2455 1830
rect 2473 1818 2476 1830
rect 2489 1818 2492 1830
rect 2503 1821 2515 1824
rect 2531 1818 2534 1830
rect 2547 1818 2550 1830
rect 2568 1818 2571 1830
rect 2584 1818 2587 1830
rect 2605 1818 2608 1830
rect 2621 1818 2624 1830
rect 2635 1821 2647 1824
rect 2663 1818 2666 1830
rect 2679 1818 2682 1830
rect 2700 1818 2703 1830
rect 2716 1818 2719 1830
rect 2737 1818 2740 1830
rect 2753 1818 2756 1830
rect 2767 1821 2779 1824
rect 2795 1818 2798 1830
rect 2811 1818 2814 1830
rect 2832 1818 2835 1830
rect 1504 1814 1537 1818
rect 1541 1814 1565 1818
rect 1569 1814 1595 1818
rect 1599 1814 1669 1818
rect 1673 1814 1697 1818
rect 1701 1814 1727 1818
rect 1731 1814 1801 1818
rect 1805 1814 1829 1818
rect 1833 1814 1859 1818
rect 1863 1814 1916 1818
rect 2449 1814 2482 1818
rect 2486 1814 2510 1818
rect 2514 1814 2540 1818
rect 2544 1814 2614 1818
rect 2618 1814 2642 1818
rect 2646 1814 2672 1818
rect 2676 1814 2746 1818
rect 2750 1814 2774 1818
rect 2778 1814 2804 1818
rect 2808 1814 2861 1818
rect 1504 1807 1513 1811
rect 1517 1807 1564 1811
rect 1568 1807 1614 1811
rect 1618 1807 1645 1811
rect 1649 1807 1696 1811
rect 1700 1807 1746 1811
rect 1750 1807 1777 1811
rect 1781 1807 1828 1811
rect 1832 1807 1878 1811
rect 1882 1807 1952 1811
rect 2449 1807 2458 1811
rect 2462 1807 2509 1811
rect 2513 1807 2559 1811
rect 2563 1807 2590 1811
rect 2594 1807 2641 1811
rect 2645 1807 2691 1811
rect 2695 1807 2722 1811
rect 2726 1807 2773 1811
rect 2777 1807 2823 1811
rect 2827 1807 2897 1811
<< m2contact >>
rect 2027 4300 2040 4304
rect 2645 4312 2658 4316
rect 2336 4300 2349 4304
rect 2691 4298 2695 4302
rect 2990 4299 2994 4314
rect 2736 4273 2740 4277
rect 2690 4259 2694 4263
rect 2705 4259 2709 4263
rect 2713 4251 2717 4255
rect 2744 4251 2748 4259
rect 2726 4237 2730 4241
rect 2998 4264 3002 4279
rect 3006 4246 3010 4259
rect 2923 4231 2927 4235
rect 2956 4231 2960 4235
rect 2990 4200 2995 4204
rect 2736 4193 2740 4197
rect 2656 4178 2660 4182
rect 2744 4177 2748 4181
rect 2726 4157 2730 4161
rect 2998 4150 3002 4154
rect 2736 4143 2740 4147
rect 2668 4129 2672 4133
rect 2683 4129 2687 4133
rect 2690 4129 2694 4133
rect 2705 4129 2709 4133
rect 2713 4121 2717 4125
rect 2744 4121 2748 4129
rect 2726 4107 2730 4111
rect 2818 4101 2822 4105
rect 2862 4102 2866 4106
rect 2990 4070 2995 4074
rect 2736 4063 2740 4067
rect 2658 4048 2662 4052
rect 2744 4047 2748 4051
rect 2726 4027 2730 4031
rect 2998 4020 3002 4024
rect 2861 3994 2867 3998
rect 2923 3994 2927 3998
rect 2873 3987 2879 3991
rect 2930 3987 2934 3991
rect 1897 3962 1901 3966
rect 2027 3962 2040 3966
rect 1987 3951 1991 3955
rect 2336 3951 2349 3955
rect 1964 3943 1970 3947
rect 2897 3943 2903 3947
rect 1952 3935 1958 3939
rect 2885 3935 2891 3939
rect 1940 3928 1946 3932
rect 2873 3928 2879 3932
rect 1928 3921 1934 3925
rect 2861 3921 2867 3925
rect 1916 3912 1922 3917
rect 2849 3913 2855 3917
rect 2990 3913 2995 3917
rect 1904 3905 1910 3909
rect 2837 3906 2843 3910
rect 2998 3906 3002 3910
rect 1976 3898 1982 3902
rect 2921 3898 2927 3902
rect 3006 3898 3010 3902
rect 2897 3836 2903 3840
rect 2909 3836 2915 3840
rect 2885 3828 2891 3832
rect 2897 3828 2903 3832
rect 2873 3820 2879 3824
rect 2885 3820 2891 3824
rect 1616 3815 1620 3819
rect 1897 3815 1901 3819
rect 2861 3812 2867 3816
rect 2873 3812 2879 3816
rect 1638 3807 1642 3811
rect 1987 3807 1991 3811
rect 2849 3804 2855 3808
rect 2861 3804 2867 3808
rect 2837 3796 2843 3800
rect 2849 3796 2855 3800
rect 1964 3763 1970 3767
rect 1997 3763 2001 3767
rect 2033 3763 2037 3767
rect 2100 3763 2104 3767
rect 2129 3763 2133 3767
rect 2165 3763 2169 3767
rect 2232 3763 2236 3767
rect 2261 3763 2265 3767
rect 2297 3763 2301 3767
rect 2364 3763 2368 3767
rect 2393 3763 2397 3767
rect 2429 3763 2433 3767
rect 2496 3763 2500 3767
rect 2909 3763 2915 3767
rect 2942 3763 2946 3767
rect 2978 3763 2982 3767
rect 3045 3763 3049 3767
rect 3074 3763 3078 3767
rect 3110 3763 3114 3767
rect 3177 3763 3181 3767
rect 3206 3763 3210 3767
rect 3242 3763 3246 3767
rect 3309 3763 3313 3767
rect 3338 3763 3342 3767
rect 3374 3763 3378 3767
rect 3441 3763 3445 3767
rect 1904 3756 1910 3760
rect 2849 3756 2855 3760
rect 1997 3749 2001 3753
rect 2047 3749 2051 3753
rect 2100 3749 2104 3753
rect 2129 3749 2133 3753
rect 2179 3749 2183 3753
rect 2232 3749 2236 3753
rect 2261 3749 2265 3753
rect 2311 3749 2315 3753
rect 2364 3749 2368 3753
rect 2393 3749 2397 3753
rect 2443 3749 2447 3753
rect 2496 3749 2500 3753
rect 2942 3749 2946 3753
rect 2992 3749 2996 3753
rect 3045 3749 3049 3753
rect 3074 3749 3078 3753
rect 3124 3749 3128 3753
rect 3177 3749 3181 3753
rect 3206 3749 3210 3753
rect 3256 3749 3260 3753
rect 3309 3749 3313 3753
rect 3338 3749 3342 3753
rect 3388 3749 3392 3753
rect 3441 3749 3445 3753
rect 2020 3738 2024 3742
rect 1645 3730 1649 3734
rect 1681 3730 1685 3734
rect 1748 3730 1752 3734
rect 1964 3730 1970 3734
rect 1991 3729 1995 3733
rect 2004 3732 2008 3738
rect 2041 3732 2045 3738
rect 2054 3734 2058 3738
rect 2078 3738 2082 3742
rect 2152 3738 2156 3742
rect 2062 3732 2066 3738
rect 2099 3732 2103 3738
rect 2115 3734 2119 3738
rect 1904 3723 1910 3727
rect 1645 3716 1649 3720
rect 1695 3716 1699 3720
rect 1748 3716 1752 3720
rect 2004 3719 2008 3723
rect 2020 3719 2024 3725
rect 2054 3725 2058 3729
rect 2041 3719 2045 3723
rect 2062 3719 2066 3723
rect 2078 3719 2082 3725
rect 2123 3729 2127 3733
rect 2136 3732 2140 3738
rect 2173 3732 2177 3738
rect 2186 3734 2190 3738
rect 2210 3738 2214 3742
rect 2284 3738 2288 3742
rect 2194 3732 2198 3738
rect 2231 3732 2235 3738
rect 2247 3734 2251 3738
rect 2099 3719 2103 3723
rect 2115 3719 2119 3723
rect 2136 3719 2140 3723
rect 2152 3719 2156 3725
rect 2186 3725 2190 3729
rect 2173 3719 2177 3723
rect 2194 3719 2198 3723
rect 2210 3719 2214 3725
rect 2255 3729 2259 3733
rect 2268 3732 2272 3738
rect 2305 3732 2309 3738
rect 2318 3734 2322 3738
rect 2342 3738 2346 3742
rect 2416 3738 2420 3742
rect 2326 3732 2330 3738
rect 2363 3732 2367 3738
rect 2379 3734 2383 3738
rect 2231 3719 2235 3723
rect 2247 3719 2251 3723
rect 2268 3719 2272 3723
rect 2284 3719 2288 3725
rect 2318 3725 2322 3729
rect 2305 3719 2309 3723
rect 2326 3719 2330 3723
rect 2342 3719 2346 3725
rect 2387 3729 2391 3733
rect 2400 3732 2404 3738
rect 2437 3732 2441 3738
rect 2450 3734 2454 3738
rect 2474 3738 2478 3742
rect 2965 3738 2969 3742
rect 2458 3732 2462 3738
rect 2495 3732 2499 3738
rect 2511 3734 2515 3738
rect 2590 3730 2594 3734
rect 2626 3730 2630 3734
rect 2693 3730 2697 3734
rect 2909 3730 2915 3734
rect 2363 3719 2367 3723
rect 2379 3719 2383 3723
rect 2400 3719 2404 3723
rect 2416 3719 2420 3725
rect 2450 3725 2454 3729
rect 2437 3719 2441 3723
rect 1668 3705 1672 3709
rect 1630 3696 1634 3700
rect 1652 3699 1656 3705
rect 1689 3699 1693 3705
rect 1702 3701 1706 3705
rect 1726 3705 1730 3709
rect 1710 3699 1714 3705
rect 1747 3699 1751 3705
rect 1763 3699 1767 3705
rect 1997 3708 2001 3712
rect 2034 3706 2038 3710
rect 2054 3706 2058 3710
rect 2098 3706 2102 3710
rect 2129 3708 2133 3712
rect 2166 3706 2170 3710
rect 2186 3706 2190 3710
rect 2230 3706 2234 3710
rect 2261 3708 2265 3712
rect 2298 3706 2302 3710
rect 2318 3706 2322 3710
rect 2362 3706 2366 3710
rect 2379 3711 2383 3715
rect 2458 3719 2462 3723
rect 2474 3719 2478 3725
rect 2936 3729 2940 3733
rect 2949 3732 2953 3738
rect 2986 3732 2990 3738
rect 2999 3734 3003 3738
rect 3023 3738 3027 3742
rect 3097 3738 3101 3742
rect 3007 3732 3011 3738
rect 3044 3732 3048 3738
rect 3060 3734 3064 3738
rect 2849 3723 2855 3727
rect 2495 3719 2499 3723
rect 2511 3719 2515 3723
rect 2393 3708 2397 3712
rect 2430 3706 2434 3710
rect 2450 3706 2454 3710
rect 2494 3706 2498 3710
rect 2511 3711 2515 3715
rect 2590 3716 2594 3720
rect 2640 3716 2644 3720
rect 2693 3716 2697 3720
rect 2949 3719 2953 3723
rect 2965 3719 2969 3725
rect 2999 3725 3003 3729
rect 2986 3719 2990 3723
rect 3007 3719 3011 3723
rect 3023 3719 3027 3725
rect 3068 3729 3072 3733
rect 3081 3732 3085 3738
rect 3118 3732 3122 3738
rect 3131 3734 3135 3738
rect 3155 3738 3159 3742
rect 3229 3738 3233 3742
rect 3139 3732 3143 3738
rect 3176 3732 3180 3738
rect 3192 3734 3196 3738
rect 3044 3719 3048 3723
rect 3060 3719 3064 3723
rect 3081 3719 3085 3723
rect 3097 3719 3101 3725
rect 3131 3725 3135 3729
rect 3118 3719 3122 3723
rect 3139 3719 3143 3723
rect 3155 3719 3159 3725
rect 3200 3729 3204 3733
rect 3213 3732 3217 3738
rect 3250 3732 3254 3738
rect 3263 3734 3267 3738
rect 3287 3738 3291 3742
rect 3361 3738 3365 3742
rect 3271 3732 3275 3738
rect 3308 3732 3312 3738
rect 3324 3734 3328 3738
rect 3176 3719 3180 3723
rect 3192 3719 3196 3723
rect 3213 3719 3217 3723
rect 3229 3719 3233 3725
rect 3263 3725 3267 3729
rect 3250 3719 3254 3723
rect 3271 3719 3275 3723
rect 3287 3719 3291 3725
rect 3332 3729 3336 3733
rect 3345 3732 3349 3738
rect 3382 3732 3386 3738
rect 3395 3734 3399 3738
rect 3419 3738 3423 3742
rect 3403 3732 3407 3738
rect 3440 3732 3444 3738
rect 3456 3734 3460 3738
rect 3308 3719 3312 3723
rect 3324 3719 3328 3723
rect 3345 3719 3349 3723
rect 3361 3719 3365 3725
rect 3395 3725 3399 3729
rect 3382 3719 3386 3723
rect 2613 3705 2617 3709
rect 1916 3699 1922 3703
rect 1652 3686 1656 3690
rect 1668 3686 1672 3692
rect 1702 3692 1706 3696
rect 1689 3686 1693 3690
rect 1710 3686 1714 3690
rect 1726 3686 1730 3692
rect 2575 3696 2579 3700
rect 2597 3699 2601 3705
rect 2634 3699 2638 3705
rect 2647 3701 2651 3705
rect 2671 3705 2675 3709
rect 2655 3699 2659 3705
rect 2692 3699 2696 3705
rect 2708 3699 2712 3705
rect 2942 3708 2946 3712
rect 2979 3706 2983 3710
rect 2999 3706 3003 3710
rect 3043 3706 3047 3710
rect 3074 3708 3078 3712
rect 3111 3706 3115 3710
rect 3131 3706 3135 3710
rect 3175 3706 3179 3710
rect 3206 3708 3210 3712
rect 3243 3706 3247 3710
rect 3263 3706 3267 3710
rect 3307 3706 3311 3710
rect 3324 3711 3328 3715
rect 3403 3719 3407 3723
rect 3419 3719 3423 3725
rect 3440 3719 3444 3723
rect 3456 3719 3460 3723
rect 3338 3708 3342 3712
rect 3375 3706 3379 3710
rect 3395 3706 3399 3710
rect 3439 3706 3443 3710
rect 3456 3711 3460 3715
rect 2861 3699 2867 3703
rect 1952 3692 1958 3696
rect 1997 3692 2001 3696
rect 2048 3692 2052 3696
rect 2098 3692 2102 3696
rect 2129 3692 2133 3696
rect 2180 3692 2184 3696
rect 2230 3692 2234 3696
rect 2261 3692 2265 3696
rect 2312 3692 2316 3696
rect 2362 3692 2366 3696
rect 2393 3692 2397 3696
rect 2444 3692 2448 3696
rect 2494 3692 2498 3696
rect 1747 3686 1751 3690
rect 1763 3686 1767 3690
rect 2597 3686 2601 3690
rect 2613 3686 2617 3692
rect 2647 3692 2651 3696
rect 2634 3686 2638 3690
rect 1645 3675 1649 3679
rect 1682 3673 1686 3677
rect 1702 3673 1706 3677
rect 1746 3673 1750 3677
rect 1904 3679 1910 3683
rect 1995 3679 1999 3683
rect 2029 3679 2033 3683
rect 2046 3679 2050 3683
rect 2102 3679 2106 3683
rect 2119 3679 2123 3683
rect 2147 3679 2151 3683
rect 2655 3686 2659 3690
rect 2671 3686 2675 3692
rect 2897 3692 2903 3696
rect 2942 3692 2946 3696
rect 2993 3692 2997 3696
rect 3043 3692 3047 3696
rect 3074 3692 3078 3696
rect 3125 3692 3129 3696
rect 3175 3692 3179 3696
rect 3206 3692 3210 3696
rect 3257 3692 3261 3696
rect 3307 3692 3311 3696
rect 3338 3692 3342 3696
rect 3389 3692 3393 3696
rect 3439 3692 3443 3696
rect 2692 3686 2696 3690
rect 2708 3686 2712 3690
rect 1940 3672 1946 3676
rect 2022 3672 2026 3676
rect 2053 3672 2057 3676
rect 2075 3672 2079 3676
rect 2140 3672 2144 3676
rect 1916 3666 1922 3670
rect 1645 3659 1649 3663
rect 1696 3659 1700 3663
rect 1746 3659 1750 3663
rect 1952 3659 1958 3663
rect 1996 3662 2000 3666
rect 2021 3665 2025 3669
rect 2028 3662 2032 3666
rect 2046 3662 2050 3666
rect 2068 3665 2072 3669
rect 2093 3665 2097 3669
rect 2103 3662 2107 3666
rect 2119 3662 2123 3666
rect 2139 3665 2143 3669
rect 2146 3662 2150 3666
rect 2210 3672 2214 3676
rect 1763 3652 1767 3656
rect 1630 3643 1634 3647
rect 1755 3645 1759 3649
rect 1779 3645 1783 3649
rect 1638 3636 1642 3640
rect 1779 3636 1783 3640
rect 2023 3646 2027 3650
rect 2043 3643 2047 3647
rect 2062 3647 2066 3651
rect 2164 3658 2168 3662
rect 2179 3658 2183 3662
rect 2081 3646 2085 3650
rect 2100 3646 2104 3650
rect 2113 3645 2117 3649
rect 2135 3646 2139 3650
rect 2143 3645 2147 3649
rect 2155 3645 2159 3649
rect 1996 3632 2000 3636
rect 2028 3632 2032 3636
rect 2046 3632 2050 3636
rect 2103 3632 2107 3636
rect 2118 3632 2122 3636
rect 2146 3632 2150 3636
rect 1645 3628 1649 3632
rect 1712 3628 1716 3632
rect 1748 3628 1752 3632
rect 1964 3628 1970 3632
rect 2010 3628 2014 3632
rect 2053 3627 2057 3631
rect 2075 3628 2082 3632
rect 2125 3627 2129 3631
rect 1904 3621 1910 3625
rect 1645 3614 1649 3618
rect 1698 3614 1702 3618
rect 1748 3614 1752 3618
rect 1928 3620 1934 3624
rect 2010 3620 2014 3624
rect 2069 3620 2073 3624
rect 2094 3620 2098 3624
rect 2125 3620 2129 3624
rect 2218 3650 2222 3658
rect 2291 3672 2295 3676
rect 2245 3658 2249 3662
rect 2260 3658 2264 3662
rect 2590 3675 2594 3679
rect 2627 3673 2631 3677
rect 2647 3673 2651 3677
rect 2691 3673 2695 3677
rect 2849 3679 2855 3683
rect 2940 3679 2944 3683
rect 2974 3679 2978 3683
rect 2991 3679 2995 3683
rect 3047 3679 3051 3683
rect 3064 3679 3068 3683
rect 3092 3679 3096 3683
rect 2885 3672 2891 3676
rect 2967 3672 2971 3676
rect 2998 3672 3002 3676
rect 3020 3672 3024 3676
rect 3085 3672 3089 3676
rect 2241 3650 2245 3654
rect 2187 3644 2191 3648
rect 2200 3636 2204 3640
rect 2299 3650 2303 3658
rect 2861 3666 2867 3670
rect 2590 3659 2594 3663
rect 2641 3659 2645 3663
rect 2691 3659 2695 3663
rect 2897 3659 2903 3663
rect 2941 3662 2945 3666
rect 2966 3665 2970 3669
rect 2973 3662 2977 3666
rect 2991 3662 2995 3666
rect 3013 3665 3017 3669
rect 3038 3665 3042 3669
rect 3048 3662 3052 3666
rect 3064 3662 3068 3666
rect 3084 3665 3088 3669
rect 3091 3662 3095 3666
rect 3155 3672 3159 3676
rect 2326 3650 2330 3654
rect 2708 3652 2712 3656
rect 2268 3644 2272 3648
rect 2575 3643 2579 3647
rect 2700 3645 2704 3649
rect 2724 3645 2728 3649
rect 2933 3645 2937 3649
rect 2281 3636 2285 3640
rect 2583 3636 2587 3640
rect 2724 3636 2728 3640
rect 2968 3646 2972 3650
rect 2988 3643 2992 3647
rect 3007 3647 3011 3651
rect 3109 3658 3113 3662
rect 3124 3658 3128 3662
rect 3026 3646 3030 3650
rect 3045 3646 3049 3650
rect 3058 3645 3062 3649
rect 3080 3646 3084 3650
rect 3088 3645 3092 3649
rect 3100 3645 3104 3649
rect 2941 3632 2945 3636
rect 2973 3632 2977 3636
rect 2991 3632 2995 3636
rect 3048 3632 3052 3636
rect 3063 3632 3067 3636
rect 3091 3632 3095 3636
rect 2590 3628 2594 3632
rect 2657 3628 2661 3632
rect 2693 3628 2697 3632
rect 2909 3628 2915 3632
rect 2955 3628 2959 3632
rect 2998 3627 3002 3631
rect 3020 3628 3027 3632
rect 3070 3627 3074 3631
rect 2849 3621 2855 3625
rect 1916 3613 1922 3617
rect 1996 3613 2000 3617
rect 2010 3613 2014 3617
rect 2028 3613 2032 3617
rect 2046 3613 2050 3617
rect 2069 3613 2073 3617
rect 2103 3613 2107 3617
rect 2118 3613 2122 3617
rect 2146 3613 2150 3617
rect 1667 3603 1671 3607
rect 1630 3597 1634 3603
rect 1646 3597 1650 3603
rect 1683 3597 1687 3603
rect 1691 3599 1695 3603
rect 1725 3603 1729 3607
rect 1928 3606 1934 3610
rect 2010 3606 2014 3610
rect 2069 3606 2073 3610
rect 2094 3606 2098 3610
rect 2125 3606 2129 3610
rect 1704 3597 1708 3603
rect 1741 3597 1745 3603
rect 2010 3598 2014 3602
rect 2053 3599 2057 3603
rect 2075 3598 2082 3602
rect 2125 3599 2129 3603
rect 1763 3594 1767 3598
rect 1996 3594 2000 3598
rect 2028 3594 2032 3598
rect 2046 3594 2050 3598
rect 2103 3594 2107 3598
rect 2118 3594 2122 3598
rect 2146 3594 2150 3598
rect 1630 3584 1634 3588
rect 1646 3584 1650 3588
rect 1691 3590 1695 3594
rect 1667 3584 1671 3590
rect 1683 3584 1687 3588
rect 1704 3584 1708 3588
rect 1725 3584 1729 3590
rect 1741 3584 1745 3588
rect 1991 3582 1995 3586
rect 1647 3571 1651 3575
rect 1691 3571 1695 3575
rect 1711 3571 1715 3575
rect 1748 3573 1752 3577
rect 2023 3580 2027 3584
rect 2043 3583 2047 3587
rect 2062 3579 2066 3583
rect 2081 3580 2085 3584
rect 2100 3580 2104 3584
rect 2113 3581 2117 3585
rect 2210 3596 2214 3600
rect 2590 3614 2594 3618
rect 2643 3614 2647 3618
rect 2693 3614 2697 3618
rect 2873 3620 2879 3624
rect 2955 3620 2959 3624
rect 3014 3620 3018 3624
rect 3039 3620 3043 3624
rect 3070 3620 3074 3624
rect 3163 3650 3167 3658
rect 3236 3672 3240 3676
rect 3190 3658 3194 3662
rect 3205 3658 3209 3662
rect 3186 3650 3190 3654
rect 3132 3644 3136 3648
rect 3145 3636 3149 3640
rect 3244 3650 3248 3658
rect 3271 3650 3275 3654
rect 3213 3644 3217 3648
rect 3226 3636 3230 3640
rect 2861 3613 2867 3617
rect 2941 3613 2945 3617
rect 2955 3613 2959 3617
rect 2973 3613 2977 3617
rect 2991 3613 2995 3617
rect 3014 3613 3018 3617
rect 3048 3613 3052 3617
rect 3063 3613 3067 3617
rect 3091 3613 3095 3617
rect 2612 3603 2616 3607
rect 2291 3596 2295 3600
rect 2575 3597 2579 3603
rect 2591 3597 2595 3603
rect 2628 3597 2632 3603
rect 2636 3599 2640 3603
rect 2670 3603 2674 3607
rect 2873 3606 2879 3610
rect 2955 3606 2959 3610
rect 3014 3606 3018 3610
rect 3039 3606 3043 3610
rect 3070 3606 3074 3610
rect 2649 3597 2653 3603
rect 2686 3597 2690 3603
rect 2955 3598 2959 3602
rect 2998 3599 3002 3603
rect 3020 3598 3027 3602
rect 3070 3599 3074 3603
rect 2708 3594 2712 3598
rect 2941 3594 2945 3598
rect 2973 3594 2977 3598
rect 2991 3594 2995 3598
rect 3048 3594 3052 3598
rect 3063 3594 3067 3598
rect 3091 3594 3095 3598
rect 2135 3580 2139 3584
rect 2143 3581 2147 3585
rect 2155 3581 2159 3585
rect 2190 3581 2194 3585
rect 2218 3580 2222 3584
rect 2270 3581 2274 3585
rect 2575 3584 2579 3588
rect 2591 3584 2595 3588
rect 2636 3590 2640 3594
rect 2612 3584 2616 3590
rect 2628 3584 2632 3588
rect 2299 3580 2303 3584
rect 2649 3584 2653 3588
rect 2670 3584 2674 3590
rect 2686 3584 2690 3588
rect 2936 3582 2940 3586
rect 1916 3564 1922 3568
rect 1996 3564 2000 3568
rect 2021 3561 2025 3565
rect 2028 3564 2032 3568
rect 2046 3564 2050 3568
rect 2068 3561 2072 3565
rect 2093 3561 2097 3565
rect 2103 3564 2107 3568
rect 2119 3564 2123 3568
rect 2139 3561 2143 3565
rect 2146 3564 2150 3568
rect 1647 3557 1651 3561
rect 1697 3557 1701 3561
rect 1748 3557 1752 3561
rect 1952 3557 1958 3561
rect 2006 3554 2010 3558
rect 2022 3554 2026 3558
rect 2053 3554 2057 3558
rect 2075 3554 2079 3558
rect 2140 3554 2144 3558
rect 2200 3560 2204 3564
rect 2592 3571 2596 3575
rect 2636 3571 2640 3575
rect 2656 3571 2660 3575
rect 2693 3573 2697 3577
rect 2968 3580 2972 3584
rect 2988 3583 2992 3587
rect 3007 3579 3011 3583
rect 3026 3580 3030 3584
rect 3045 3580 3049 3584
rect 3058 3581 3062 3585
rect 3155 3596 3159 3600
rect 3236 3596 3240 3600
rect 3080 3580 3084 3584
rect 3088 3581 3092 3585
rect 3100 3581 3104 3585
rect 3135 3581 3139 3585
rect 3163 3580 3167 3584
rect 3215 3581 3219 3585
rect 3244 3580 3248 3584
rect 2861 3564 2867 3568
rect 2941 3564 2945 3568
rect 2281 3560 2285 3564
rect 2966 3561 2970 3565
rect 2973 3564 2977 3568
rect 2991 3564 2995 3568
rect 3013 3561 3017 3565
rect 3038 3561 3042 3565
rect 3048 3564 3052 3568
rect 3064 3564 3068 3568
rect 3084 3561 3088 3565
rect 3091 3564 3095 3568
rect 2592 3557 2596 3561
rect 2642 3557 2646 3561
rect 2693 3557 2697 3561
rect 2897 3557 2903 3561
rect 2951 3554 2955 3558
rect 2967 3554 2971 3558
rect 2998 3554 3002 3558
rect 3020 3554 3024 3558
rect 3085 3554 3089 3558
rect 3145 3560 3149 3564
rect 3226 3560 3230 3564
rect 1904 3547 1910 3551
rect 1995 3547 1999 3551
rect 2029 3547 2033 3551
rect 2046 3547 2050 3551
rect 2102 3547 2106 3551
rect 2119 3547 2123 3551
rect 2147 3547 2151 3551
rect 2849 3547 2855 3551
rect 2940 3547 2944 3551
rect 2974 3547 2978 3551
rect 2991 3547 2995 3551
rect 3047 3547 3051 3551
rect 3064 3547 3068 3551
rect 3092 3547 3096 3551
rect 1940 3540 1946 3544
rect 2006 3540 2010 3544
rect 2022 3540 2026 3544
rect 2053 3540 2057 3544
rect 2075 3540 2079 3544
rect 2140 3540 2144 3544
rect 2210 3540 2214 3544
rect 1996 3530 2000 3534
rect 2021 3533 2025 3537
rect 2028 3530 2032 3534
rect 2046 3530 2050 3534
rect 2068 3533 2072 3537
rect 2093 3533 2097 3537
rect 2103 3530 2107 3534
rect 2119 3530 2123 3534
rect 2139 3533 2143 3537
rect 2146 3530 2150 3534
rect 1990 3513 1994 3517
rect 2023 3514 2027 3518
rect 2043 3511 2047 3515
rect 2062 3515 2066 3519
rect 2081 3514 2085 3518
rect 2100 3514 2104 3518
rect 2113 3513 2117 3517
rect 2135 3514 2139 3518
rect 2143 3513 2147 3517
rect 2155 3513 2159 3517
rect 2218 3518 2222 3526
rect 2315 3540 2319 3544
rect 2269 3526 2273 3530
rect 2284 3526 2288 3530
rect 2885 3540 2891 3544
rect 2951 3540 2955 3544
rect 2967 3540 2971 3544
rect 2998 3540 3002 3544
rect 3020 3540 3024 3544
rect 3085 3540 3089 3544
rect 3155 3540 3159 3544
rect 2187 3512 2191 3516
rect 2241 3517 2245 3521
rect 1996 3500 2000 3504
rect 2028 3500 2032 3504
rect 2046 3500 2050 3504
rect 2103 3500 2107 3504
rect 2118 3500 2122 3504
rect 2146 3500 2150 3504
rect 2010 3496 2014 3500
rect 2053 3495 2057 3499
rect 2075 3496 2082 3500
rect 2125 3495 2129 3499
rect 1928 3488 1934 3492
rect 2010 3488 2014 3492
rect 2069 3488 2073 3492
rect 2094 3488 2098 3492
rect 2125 3488 2129 3492
rect 2200 3504 2204 3508
rect 2323 3518 2327 3526
rect 2941 3530 2945 3534
rect 2966 3533 2970 3537
rect 2973 3530 2977 3534
rect 2991 3530 2995 3534
rect 3013 3533 3017 3537
rect 3038 3533 3042 3537
rect 3048 3530 3052 3534
rect 3064 3530 3068 3534
rect 3084 3533 3088 3537
rect 3091 3530 3095 3534
rect 2344 3518 2348 3522
rect 2292 3512 2296 3516
rect 2935 3513 2939 3517
rect 2305 3504 2309 3508
rect 2968 3514 2972 3518
rect 2988 3511 2992 3515
rect 3007 3515 3011 3519
rect 3026 3514 3030 3518
rect 3045 3514 3049 3518
rect 3058 3513 3062 3517
rect 3080 3514 3084 3518
rect 3088 3513 3092 3517
rect 3100 3513 3104 3517
rect 3163 3518 3167 3526
rect 3260 3540 3264 3544
rect 3214 3526 3218 3530
rect 3229 3526 3233 3530
rect 3132 3512 3136 3516
rect 3186 3517 3190 3521
rect 2941 3500 2945 3504
rect 2973 3500 2977 3504
rect 2991 3500 2995 3504
rect 3048 3500 3052 3504
rect 3063 3500 3067 3504
rect 3091 3500 3095 3504
rect 2955 3496 2959 3500
rect 2998 3495 3002 3499
rect 3020 3496 3027 3500
rect 3070 3495 3074 3499
rect 2873 3488 2879 3492
rect 2955 3488 2959 3492
rect 3014 3488 3018 3492
rect 3039 3488 3043 3492
rect 3070 3488 3074 3492
rect 3145 3504 3149 3508
rect 3268 3518 3272 3526
rect 3289 3518 3293 3522
rect 3237 3512 3241 3516
rect 3250 3504 3254 3508
rect 1916 3481 1922 3485
rect 1996 3481 2000 3485
rect 2010 3481 2014 3485
rect 2028 3481 2032 3485
rect 2046 3481 2050 3485
rect 2069 3481 2073 3485
rect 2103 3481 2107 3485
rect 2118 3481 2122 3485
rect 2146 3481 2150 3485
rect 2861 3481 2867 3485
rect 2941 3481 2945 3485
rect 2955 3481 2959 3485
rect 2973 3481 2977 3485
rect 2991 3481 2995 3485
rect 3014 3481 3018 3485
rect 3048 3481 3052 3485
rect 3063 3481 3067 3485
rect 3091 3481 3095 3485
rect 1928 3474 1934 3478
rect 2010 3474 2014 3478
rect 2069 3474 2073 3478
rect 2094 3474 2098 3478
rect 2125 3474 2129 3478
rect 2010 3466 2014 3470
rect 2053 3467 2057 3471
rect 2075 3466 2082 3470
rect 2125 3467 2129 3471
rect 1996 3462 2000 3466
rect 2028 3462 2032 3466
rect 2046 3462 2050 3466
rect 2103 3462 2107 3466
rect 2118 3462 2122 3466
rect 2146 3462 2150 3466
rect 2210 3465 2214 3469
rect 2873 3474 2879 3478
rect 2955 3474 2959 3478
rect 3014 3474 3018 3478
rect 3039 3474 3043 3478
rect 3070 3474 3074 3478
rect 2315 3465 2319 3469
rect 2955 3466 2959 3470
rect 2998 3467 3002 3471
rect 3020 3466 3027 3470
rect 3070 3467 3074 3471
rect 2941 3462 2945 3466
rect 2973 3462 2977 3466
rect 2991 3462 2995 3466
rect 3048 3462 3052 3466
rect 3063 3462 3067 3466
rect 3091 3462 3095 3466
rect 3155 3465 3159 3469
rect 3260 3465 3264 3469
rect 1991 3450 1995 3454
rect 2023 3448 2027 3452
rect 2043 3451 2047 3455
rect 2062 3447 2066 3451
rect 2081 3448 2085 3452
rect 2100 3448 2104 3452
rect 2113 3449 2117 3453
rect 2135 3448 2139 3452
rect 2143 3449 2147 3453
rect 2155 3449 2159 3453
rect 2189 3450 2193 3454
rect 2218 3449 2222 3453
rect 2295 3450 2299 3454
rect 2323 3449 2327 3453
rect 2936 3450 2940 3454
rect 1996 3432 2000 3436
rect 2021 3429 2025 3433
rect 2028 3432 2032 3436
rect 2046 3432 2050 3436
rect 2068 3429 2072 3433
rect 2093 3429 2097 3433
rect 2103 3432 2107 3436
rect 2119 3432 2123 3436
rect 2139 3429 2143 3433
rect 2146 3432 2150 3436
rect 1940 3422 1946 3426
rect 2022 3422 2026 3426
rect 2053 3422 2057 3426
rect 2075 3422 2079 3426
rect 2140 3422 2144 3426
rect 2200 3429 2204 3433
rect 2968 3448 2972 3452
rect 2988 3451 2992 3455
rect 3007 3447 3011 3451
rect 3026 3448 3030 3452
rect 3045 3448 3049 3452
rect 3058 3449 3062 3453
rect 3080 3448 3084 3452
rect 3088 3449 3092 3453
rect 3100 3449 3104 3453
rect 3134 3450 3138 3454
rect 3163 3449 3167 3453
rect 3240 3450 3244 3454
rect 3268 3449 3272 3453
rect 2305 3429 2309 3433
rect 2941 3432 2945 3436
rect 2966 3429 2970 3433
rect 2973 3432 2977 3436
rect 2991 3432 2995 3436
rect 3013 3429 3017 3433
rect 3038 3429 3042 3433
rect 3048 3432 3052 3436
rect 3064 3432 3068 3436
rect 3084 3429 3088 3433
rect 3091 3432 3095 3436
rect 2885 3422 2891 3426
rect 2967 3422 2971 3426
rect 2998 3422 3002 3426
rect 3020 3422 3024 3426
rect 3085 3422 3089 3426
rect 3145 3429 3149 3433
rect 3250 3429 3254 3433
rect 1904 3415 1910 3419
rect 1995 3415 1999 3419
rect 2029 3415 2033 3419
rect 2046 3415 2050 3419
rect 2102 3415 2106 3419
rect 2119 3415 2123 3419
rect 2147 3415 2151 3419
rect 2849 3415 2855 3419
rect 2940 3415 2944 3419
rect 2974 3415 2978 3419
rect 2991 3415 2995 3419
rect 3047 3415 3051 3419
rect 3064 3415 3068 3419
rect 3092 3415 3096 3419
rect 1940 3408 1946 3412
rect 2022 3408 2026 3412
rect 2053 3408 2057 3412
rect 2075 3408 2079 3412
rect 2140 3408 2144 3412
rect 2210 3408 2214 3412
rect 1996 3398 2000 3402
rect 2021 3401 2025 3405
rect 2028 3398 2032 3402
rect 2046 3398 2050 3402
rect 2068 3401 2072 3405
rect 2093 3401 2097 3405
rect 2103 3398 2107 3402
rect 2119 3398 2123 3402
rect 2139 3401 2143 3405
rect 2146 3398 2150 3402
rect 1990 3381 1994 3385
rect 2023 3382 2027 3386
rect 2043 3379 2047 3383
rect 2062 3383 2066 3387
rect 2081 3382 2085 3386
rect 2100 3382 2104 3386
rect 2113 3381 2117 3385
rect 2135 3382 2139 3386
rect 2143 3381 2147 3385
rect 2155 3381 2159 3385
rect 2218 3386 2222 3394
rect 2291 3408 2295 3412
rect 2245 3394 2249 3398
rect 2260 3394 2264 3398
rect 2241 3386 2245 3390
rect 2187 3380 2191 3384
rect 1996 3368 2000 3372
rect 2028 3368 2032 3372
rect 2046 3368 2050 3372
rect 2103 3368 2107 3372
rect 2118 3368 2122 3372
rect 2146 3368 2150 3372
rect 2010 3364 2014 3368
rect 2053 3363 2057 3367
rect 2075 3364 2082 3368
rect 2125 3363 2129 3367
rect 1928 3356 1934 3360
rect 2010 3356 2014 3360
rect 2069 3356 2073 3360
rect 2094 3356 2098 3360
rect 2125 3356 2129 3360
rect 2200 3372 2204 3376
rect 2299 3386 2303 3394
rect 2381 3408 2385 3412
rect 2335 3394 2339 3398
rect 2350 3394 2354 3398
rect 2885 3408 2891 3412
rect 2967 3408 2971 3412
rect 2998 3408 3002 3412
rect 3020 3408 3024 3412
rect 3085 3408 3089 3412
rect 3155 3408 3159 3412
rect 2323 3386 2327 3390
rect 2268 3380 2272 3384
rect 2357 3388 2361 3392
rect 2389 3386 2393 3394
rect 2941 3398 2945 3402
rect 2966 3401 2970 3405
rect 2973 3398 2977 3402
rect 2991 3398 2995 3402
rect 3013 3401 3017 3405
rect 3038 3401 3042 3405
rect 3048 3398 3052 3402
rect 3064 3398 3068 3402
rect 3084 3401 3088 3405
rect 3091 3398 3095 3402
rect 2281 3372 2285 3376
rect 2424 3385 2428 3389
rect 2935 3381 2939 3385
rect 2371 3372 2375 3376
rect 2968 3382 2972 3386
rect 2988 3379 2992 3383
rect 3007 3383 3011 3387
rect 3026 3382 3030 3386
rect 3045 3382 3049 3386
rect 3058 3381 3062 3385
rect 3080 3382 3084 3386
rect 3088 3381 3092 3385
rect 3100 3381 3104 3385
rect 3163 3386 3167 3394
rect 3236 3408 3240 3412
rect 3190 3394 3194 3398
rect 3205 3394 3209 3398
rect 3186 3386 3190 3390
rect 3132 3380 3136 3384
rect 2941 3368 2945 3372
rect 2973 3368 2977 3372
rect 2991 3368 2995 3372
rect 3048 3368 3052 3372
rect 3063 3368 3067 3372
rect 3091 3368 3095 3372
rect 2955 3364 2959 3368
rect 2998 3363 3002 3367
rect 3020 3364 3027 3368
rect 3070 3363 3074 3367
rect 2873 3356 2879 3360
rect 2955 3356 2959 3360
rect 3014 3356 3018 3360
rect 3039 3356 3043 3360
rect 3070 3356 3074 3360
rect 3145 3372 3149 3376
rect 3244 3386 3248 3394
rect 3326 3408 3330 3412
rect 3280 3394 3284 3398
rect 3295 3394 3299 3398
rect 3268 3386 3272 3390
rect 3213 3380 3217 3384
rect 3302 3388 3306 3392
rect 3334 3386 3338 3394
rect 3226 3372 3230 3376
rect 3369 3385 3373 3389
rect 3316 3372 3320 3376
rect 1916 3349 1922 3353
rect 1996 3349 2000 3353
rect 2010 3349 2014 3353
rect 2028 3349 2032 3353
rect 2046 3349 2050 3353
rect 2069 3349 2073 3353
rect 2103 3349 2107 3353
rect 2118 3349 2122 3353
rect 2146 3349 2150 3353
rect 2861 3349 2867 3353
rect 2941 3349 2945 3353
rect 2955 3349 2959 3353
rect 2973 3349 2977 3353
rect 2991 3349 2995 3353
rect 3014 3349 3018 3353
rect 3048 3349 3052 3353
rect 3063 3349 3067 3353
rect 3091 3349 3095 3353
rect 1928 3342 1934 3346
rect 2010 3342 2014 3346
rect 2069 3342 2073 3346
rect 2094 3342 2098 3346
rect 2125 3342 2129 3346
rect 2010 3334 2014 3338
rect 2053 3335 2057 3339
rect 2075 3334 2082 3338
rect 2125 3335 2129 3339
rect 1996 3330 2000 3334
rect 2028 3330 2032 3334
rect 2046 3330 2050 3334
rect 2103 3330 2107 3334
rect 2118 3330 2122 3334
rect 2146 3330 2150 3334
rect 1991 3318 1995 3322
rect 2023 3316 2027 3320
rect 2043 3319 2047 3323
rect 2062 3315 2066 3319
rect 2081 3316 2085 3320
rect 2100 3316 2104 3320
rect 2113 3317 2117 3321
rect 2210 3330 2214 3334
rect 2291 3330 2295 3334
rect 2873 3342 2879 3346
rect 2955 3342 2959 3346
rect 3014 3342 3018 3346
rect 3039 3342 3043 3346
rect 3070 3342 3074 3346
rect 2955 3334 2959 3338
rect 2998 3335 3002 3339
rect 3020 3334 3027 3338
rect 3070 3335 3074 3339
rect 2381 3330 2385 3334
rect 2941 3330 2945 3334
rect 2973 3330 2977 3334
rect 2991 3330 2995 3334
rect 3048 3330 3052 3334
rect 3063 3330 3067 3334
rect 3091 3330 3095 3334
rect 2135 3316 2139 3320
rect 2143 3317 2147 3321
rect 2155 3317 2159 3321
rect 2190 3315 2194 3319
rect 2218 3314 2222 3318
rect 2270 3315 2274 3319
rect 2299 3314 2303 3318
rect 2354 3315 2358 3319
rect 2936 3318 2940 3322
rect 2389 3314 2393 3318
rect 1996 3300 2000 3304
rect 2021 3297 2025 3301
rect 2028 3300 2032 3304
rect 2046 3300 2050 3304
rect 2068 3297 2072 3301
rect 2093 3297 2097 3301
rect 2103 3300 2107 3304
rect 2119 3300 2123 3304
rect 2139 3297 2143 3301
rect 2146 3300 2150 3304
rect 2968 3316 2972 3320
rect 2988 3319 2992 3323
rect 3007 3315 3011 3319
rect 3026 3316 3030 3320
rect 3045 3316 3049 3320
rect 3058 3317 3062 3321
rect 3155 3330 3159 3334
rect 3236 3330 3240 3334
rect 3326 3330 3330 3334
rect 3080 3316 3084 3320
rect 3088 3317 3092 3321
rect 3100 3317 3104 3321
rect 3135 3315 3139 3319
rect 3163 3314 3167 3318
rect 3215 3315 3219 3319
rect 3244 3314 3248 3318
rect 3299 3315 3303 3319
rect 3334 3314 3338 3318
rect 1940 3290 1946 3294
rect 2022 3290 2026 3294
rect 2053 3290 2057 3294
rect 2075 3290 2079 3294
rect 2140 3290 2144 3294
rect 2200 3294 2204 3298
rect 2281 3294 2285 3298
rect 2941 3300 2945 3304
rect 2371 3294 2375 3298
rect 2966 3297 2970 3301
rect 2973 3300 2977 3304
rect 2991 3300 2995 3304
rect 3013 3297 3017 3301
rect 3038 3297 3042 3301
rect 3048 3300 3052 3304
rect 3064 3300 3068 3304
rect 3084 3297 3088 3301
rect 3091 3300 3095 3304
rect 2885 3290 2891 3294
rect 2967 3290 2971 3294
rect 2998 3290 3002 3294
rect 3020 3290 3024 3294
rect 3085 3290 3089 3294
rect 3145 3294 3149 3298
rect 3226 3294 3230 3298
rect 3316 3294 3320 3298
rect 1904 3283 1910 3287
rect 1995 3283 1999 3287
rect 2029 3283 2033 3287
rect 2046 3283 2050 3287
rect 2102 3283 2106 3287
rect 2119 3283 2123 3287
rect 2147 3283 2151 3287
rect 2849 3283 2855 3287
rect 2940 3283 2944 3287
rect 2974 3283 2978 3287
rect 2991 3283 2995 3287
rect 3047 3283 3051 3287
rect 3064 3283 3068 3287
rect 3092 3283 3096 3287
rect 1940 3276 1946 3280
rect 2022 3276 2026 3280
rect 2053 3276 2057 3280
rect 2075 3276 2079 3280
rect 2140 3276 2144 3280
rect 2210 3276 2214 3280
rect 1996 3266 2000 3270
rect 2021 3269 2025 3273
rect 2028 3266 2032 3270
rect 2046 3266 2050 3270
rect 2068 3269 2072 3273
rect 2093 3269 2097 3273
rect 2103 3266 2107 3270
rect 2119 3266 2123 3270
rect 2139 3269 2143 3273
rect 2146 3266 2150 3270
rect 1990 3249 1994 3253
rect 2023 3250 2027 3254
rect 2043 3247 2047 3251
rect 2062 3251 2066 3255
rect 2885 3276 2891 3280
rect 2967 3276 2971 3280
rect 2998 3276 3002 3280
rect 3020 3276 3024 3280
rect 3085 3276 3089 3280
rect 3155 3276 3159 3280
rect 2081 3250 2085 3254
rect 2100 3250 2104 3254
rect 2113 3249 2117 3253
rect 2135 3250 2139 3254
rect 2143 3249 2147 3253
rect 2155 3249 2159 3253
rect 2218 3254 2222 3262
rect 2941 3266 2945 3270
rect 2966 3269 2970 3273
rect 2973 3266 2977 3270
rect 2991 3266 2995 3270
rect 3013 3269 3017 3273
rect 3038 3269 3042 3273
rect 3048 3266 3052 3270
rect 3064 3266 3068 3270
rect 3084 3269 3088 3273
rect 3091 3266 3095 3270
rect 2187 3248 2191 3252
rect 2241 3253 2245 3257
rect 2935 3249 2939 3253
rect 1491 3235 1495 3239
rect 1616 3235 1620 3239
rect 1996 3236 2000 3240
rect 2028 3236 2032 3240
rect 2046 3236 2050 3240
rect 2103 3236 2107 3240
rect 2118 3236 2122 3240
rect 2146 3236 2150 3240
rect 2010 3232 2014 3236
rect 1513 3228 1517 3232
rect 1549 3228 1553 3232
rect 1616 3228 1620 3232
rect 1645 3228 1649 3232
rect 1681 3228 1685 3232
rect 1748 3228 1752 3232
rect 1777 3228 1781 3232
rect 1813 3228 1817 3232
rect 1880 3228 1884 3232
rect 1964 3228 1970 3232
rect 2053 3231 2057 3235
rect 2075 3232 2082 3236
rect 2125 3231 2129 3235
rect 1904 3221 1910 3225
rect 2010 3224 2014 3228
rect 2019 3224 2023 3228
rect 2069 3224 2073 3228
rect 2094 3224 2098 3228
rect 2125 3224 2129 3228
rect 2200 3240 2204 3244
rect 2968 3250 2972 3254
rect 2988 3247 2992 3251
rect 3007 3251 3011 3255
rect 3026 3250 3030 3254
rect 3045 3250 3049 3254
rect 3058 3249 3062 3253
rect 3080 3250 3084 3254
rect 3088 3249 3092 3253
rect 3100 3249 3104 3253
rect 3163 3254 3167 3262
rect 3132 3248 3136 3252
rect 3186 3253 3190 3257
rect 2941 3236 2945 3240
rect 2973 3236 2977 3240
rect 2991 3236 2995 3240
rect 3048 3236 3052 3240
rect 3063 3236 3067 3240
rect 3091 3236 3095 3240
rect 2955 3232 2959 3236
rect 2458 3228 2462 3232
rect 2494 3228 2498 3232
rect 2561 3228 2565 3232
rect 2590 3228 2594 3232
rect 2626 3228 2630 3232
rect 2693 3228 2697 3232
rect 2722 3228 2726 3232
rect 2758 3228 2762 3232
rect 2825 3228 2829 3232
rect 2909 3228 2915 3232
rect 2998 3231 3002 3235
rect 3020 3232 3027 3236
rect 3070 3231 3074 3235
rect 2849 3221 2855 3225
rect 2955 3224 2959 3228
rect 2964 3224 2968 3228
rect 3014 3224 3018 3228
rect 3039 3224 3043 3228
rect 3070 3224 3074 3228
rect 3145 3240 3149 3244
rect 1513 3214 1517 3218
rect 1563 3214 1567 3218
rect 1616 3214 1620 3218
rect 1645 3214 1649 3218
rect 1695 3214 1699 3218
rect 1748 3214 1752 3218
rect 1777 3214 1781 3218
rect 1827 3214 1831 3218
rect 1880 3214 1884 3218
rect 1916 3217 1922 3221
rect 1996 3217 2000 3221
rect 2010 3217 2014 3221
rect 2028 3217 2032 3221
rect 2046 3217 2050 3221
rect 2069 3217 2073 3221
rect 2103 3217 2107 3221
rect 2118 3217 2122 3221
rect 2146 3217 2150 3221
rect 2271 3217 2275 3221
rect 2289 3217 2293 3221
rect 2307 3217 2311 3221
rect 2330 3217 2334 3221
rect 2364 3217 2368 3221
rect 2379 3217 2383 3221
rect 2407 3217 2411 3221
rect 1536 3203 1540 3207
rect 1507 3194 1511 3198
rect 1520 3197 1524 3203
rect 1557 3197 1561 3203
rect 1570 3199 1574 3203
rect 1594 3203 1598 3207
rect 1668 3203 1672 3207
rect 1578 3197 1582 3203
rect 1615 3197 1619 3203
rect 1631 3197 1635 3203
rect 1652 3197 1656 3203
rect 1689 3197 1693 3203
rect 1702 3199 1706 3203
rect 1726 3203 1730 3207
rect 1800 3203 1804 3207
rect 1710 3197 1714 3203
rect 1747 3197 1751 3203
rect 1763 3197 1767 3203
rect 1784 3197 1788 3203
rect 1821 3197 1825 3203
rect 1834 3199 1838 3203
rect 1858 3203 1862 3207
rect 1928 3210 1934 3214
rect 2010 3210 2014 3214
rect 2019 3210 2023 3214
rect 2069 3210 2073 3214
rect 2094 3210 2098 3214
rect 2125 3210 2129 3214
rect 1842 3197 1846 3203
rect 1879 3197 1883 3203
rect 1895 3199 1899 3203
rect 2010 3202 2014 3206
rect 2053 3203 2057 3207
rect 2075 3202 2082 3206
rect 2125 3203 2129 3207
rect 1996 3198 2000 3202
rect 2028 3198 2032 3202
rect 2046 3198 2050 3202
rect 2103 3198 2107 3202
rect 2118 3198 2122 3202
rect 2146 3198 2150 3202
rect 1520 3184 1524 3188
rect 1536 3184 1540 3190
rect 1570 3190 1574 3194
rect 1557 3184 1561 3188
rect 1578 3184 1582 3188
rect 1594 3184 1598 3190
rect 1615 3184 1619 3188
rect 1631 3184 1635 3188
rect 1652 3184 1656 3188
rect 1668 3184 1672 3190
rect 1702 3190 1706 3194
rect 1689 3184 1693 3188
rect 1710 3184 1714 3188
rect 1726 3184 1730 3190
rect 1747 3184 1751 3188
rect 1763 3184 1767 3188
rect 1784 3184 1788 3188
rect 1800 3184 1804 3190
rect 1834 3190 1838 3194
rect 1821 3184 1825 3188
rect 1842 3184 1846 3188
rect 1858 3184 1862 3190
rect 1879 3184 1883 3188
rect 1895 3184 1899 3188
rect 1991 3186 1995 3190
rect 1513 3173 1517 3177
rect 1550 3171 1554 3175
rect 1570 3171 1574 3175
rect 1614 3171 1618 3175
rect 1645 3173 1649 3177
rect 1682 3171 1686 3175
rect 1702 3171 1706 3175
rect 1746 3171 1750 3175
rect 1777 3173 1781 3177
rect 1814 3171 1818 3175
rect 1834 3171 1838 3175
rect 1878 3171 1882 3175
rect 2023 3184 2027 3188
rect 2043 3187 2047 3191
rect 2062 3183 2066 3187
rect 2081 3184 2085 3188
rect 2100 3184 2104 3188
rect 2113 3185 2117 3189
rect 2249 3210 2253 3214
rect 2271 3210 2275 3214
rect 2330 3210 2334 3214
rect 2355 3210 2359 3214
rect 2386 3210 2390 3214
rect 2458 3214 2462 3218
rect 2508 3214 2512 3218
rect 2561 3214 2565 3218
rect 2590 3214 2594 3218
rect 2640 3214 2644 3218
rect 2693 3214 2697 3218
rect 2722 3214 2726 3218
rect 2772 3214 2776 3218
rect 2825 3214 2829 3218
rect 2861 3217 2867 3221
rect 2941 3217 2945 3221
rect 2955 3217 2959 3221
rect 2973 3217 2977 3221
rect 2991 3217 2995 3221
rect 3014 3217 3018 3221
rect 3048 3217 3052 3221
rect 3063 3217 3067 3221
rect 3091 3217 3095 3221
rect 3216 3217 3220 3221
rect 3234 3217 3238 3221
rect 3252 3217 3256 3221
rect 3275 3217 3279 3221
rect 3309 3217 3313 3221
rect 3324 3217 3328 3221
rect 3352 3217 3356 3221
rect 2271 3202 2275 3206
rect 2314 3203 2318 3207
rect 2336 3202 2343 3206
rect 2386 3203 2390 3207
rect 2481 3203 2485 3207
rect 2289 3198 2293 3202
rect 2307 3198 2311 3202
rect 2364 3198 2368 3202
rect 2379 3198 2383 3202
rect 2407 3198 2411 3202
rect 2210 3194 2214 3198
rect 2135 3184 2139 3188
rect 2143 3185 2147 3189
rect 2155 3185 2159 3189
rect 2189 3179 2193 3183
rect 2229 3185 2233 3189
rect 2218 3178 2222 3182
rect 1996 3168 2000 3172
rect 1916 3164 1922 3168
rect 2021 3165 2025 3169
rect 2028 3168 2032 3172
rect 2046 3168 2050 3172
rect 2068 3165 2072 3169
rect 2093 3165 2097 3169
rect 2103 3168 2107 3172
rect 2119 3168 2123 3172
rect 2139 3165 2143 3169
rect 2146 3168 2150 3172
rect 2284 3184 2288 3188
rect 2304 3187 2308 3191
rect 2323 3183 2327 3187
rect 2452 3194 2456 3198
rect 2465 3197 2469 3203
rect 2502 3197 2506 3203
rect 2515 3199 2519 3203
rect 2539 3203 2543 3207
rect 2613 3203 2617 3207
rect 2523 3197 2527 3203
rect 2560 3197 2564 3203
rect 2576 3197 2580 3203
rect 2597 3197 2601 3203
rect 2634 3197 2638 3203
rect 2647 3199 2651 3203
rect 2671 3203 2675 3207
rect 2745 3203 2749 3207
rect 2655 3197 2659 3203
rect 2692 3197 2696 3203
rect 2708 3197 2712 3203
rect 2729 3197 2733 3203
rect 2766 3197 2770 3203
rect 2779 3199 2783 3203
rect 2803 3203 2807 3207
rect 2873 3210 2879 3214
rect 2955 3210 2959 3214
rect 2964 3210 2968 3214
rect 3014 3210 3018 3214
rect 3039 3210 3043 3214
rect 3070 3210 3074 3214
rect 2787 3197 2791 3203
rect 2824 3197 2828 3203
rect 2840 3199 2844 3203
rect 2955 3202 2959 3206
rect 2998 3203 3002 3207
rect 3020 3202 3027 3206
rect 3070 3203 3074 3207
rect 2941 3198 2945 3202
rect 2973 3198 2977 3202
rect 2991 3198 2995 3202
rect 3048 3198 3052 3202
rect 3063 3198 3067 3202
rect 3091 3198 3095 3202
rect 2342 3184 2346 3188
rect 2361 3184 2365 3188
rect 2374 3185 2378 3189
rect 2396 3184 2400 3188
rect 2404 3185 2408 3189
rect 2416 3185 2420 3189
rect 2465 3184 2469 3188
rect 2481 3184 2485 3190
rect 2515 3190 2519 3194
rect 2502 3184 2506 3188
rect 2523 3184 2527 3188
rect 2539 3184 2543 3190
rect 2560 3184 2564 3188
rect 2576 3184 2580 3188
rect 2597 3184 2601 3188
rect 2613 3184 2617 3190
rect 2647 3190 2651 3194
rect 2634 3184 2638 3188
rect 2655 3184 2659 3188
rect 2671 3184 2675 3190
rect 2692 3184 2696 3188
rect 2708 3184 2712 3188
rect 2729 3184 2733 3188
rect 2745 3184 2749 3190
rect 2779 3190 2783 3194
rect 2766 3184 2770 3188
rect 2787 3184 2791 3188
rect 2803 3184 2807 3190
rect 2824 3184 2828 3188
rect 2840 3184 2844 3188
rect 2936 3186 2940 3190
rect 2230 3168 2234 3172
rect 2256 3168 2260 3172
rect 1513 3157 1517 3161
rect 1564 3157 1568 3161
rect 1614 3157 1618 3161
rect 1645 3157 1649 3161
rect 1696 3157 1700 3161
rect 1746 3157 1750 3161
rect 1777 3157 1781 3161
rect 1828 3157 1832 3161
rect 1878 3157 1882 3161
rect 1952 3158 1958 3162
rect 2004 3158 2008 3162
rect 2022 3158 2026 3162
rect 2053 3158 2057 3162
rect 2075 3158 2079 3162
rect 2140 3158 2144 3162
rect 2282 3165 2286 3169
rect 2289 3168 2293 3172
rect 2307 3168 2311 3172
rect 2329 3165 2333 3169
rect 2354 3165 2358 3169
rect 2364 3168 2368 3172
rect 2380 3168 2384 3172
rect 2400 3165 2404 3169
rect 2407 3168 2411 3172
rect 2458 3173 2462 3177
rect 2495 3171 2499 3175
rect 2515 3171 2519 3175
rect 2559 3171 2563 3175
rect 2590 3173 2594 3177
rect 2627 3171 2631 3175
rect 2647 3171 2651 3175
rect 2691 3171 2695 3175
rect 2722 3173 2726 3177
rect 2759 3171 2763 3175
rect 2779 3171 2783 3175
rect 2823 3171 2827 3175
rect 2968 3184 2972 3188
rect 2988 3187 2992 3191
rect 3007 3183 3011 3187
rect 3026 3184 3030 3188
rect 3045 3184 3049 3188
rect 3058 3185 3062 3189
rect 3194 3210 3198 3214
rect 3216 3210 3220 3214
rect 3275 3210 3279 3214
rect 3300 3210 3304 3214
rect 3331 3210 3335 3214
rect 3216 3202 3220 3206
rect 3259 3203 3263 3207
rect 3281 3202 3288 3206
rect 3331 3203 3335 3207
rect 3234 3198 3238 3202
rect 3252 3198 3256 3202
rect 3309 3198 3313 3202
rect 3324 3198 3328 3202
rect 3352 3198 3356 3202
rect 3155 3194 3159 3198
rect 3080 3184 3084 3188
rect 3088 3185 3092 3189
rect 3100 3185 3104 3189
rect 3134 3179 3138 3183
rect 3174 3185 3178 3189
rect 3163 3178 3167 3182
rect 2941 3168 2945 3172
rect 2861 3164 2867 3168
rect 2966 3165 2970 3169
rect 2973 3168 2977 3172
rect 2991 3168 2995 3172
rect 3013 3165 3017 3169
rect 3038 3165 3042 3169
rect 3048 3168 3052 3172
rect 3064 3168 3068 3172
rect 3084 3165 3088 3169
rect 3091 3168 3095 3172
rect 3229 3184 3233 3188
rect 3249 3187 3253 3191
rect 3268 3183 3272 3187
rect 3287 3184 3291 3188
rect 3306 3184 3310 3188
rect 3319 3185 3323 3189
rect 3341 3184 3345 3188
rect 3349 3185 3353 3189
rect 3361 3185 3365 3189
rect 3175 3168 3179 3172
rect 3201 3168 3205 3172
rect 2200 3158 2204 3162
rect 2239 3158 2243 3162
rect 2283 3158 2287 3162
rect 2314 3158 2318 3162
rect 2336 3158 2340 3162
rect 2401 3158 2405 3162
rect 2458 3157 2462 3161
rect 2509 3157 2513 3161
rect 2559 3157 2563 3161
rect 2590 3157 2594 3161
rect 2641 3157 2645 3161
rect 2691 3157 2695 3161
rect 2722 3157 2726 3161
rect 2773 3157 2777 3161
rect 2823 3157 2827 3161
rect 2897 3158 2903 3162
rect 2949 3158 2953 3162
rect 2967 3158 2971 3162
rect 2998 3158 3002 3162
rect 3020 3158 3024 3162
rect 3085 3158 3089 3162
rect 3227 3165 3231 3169
rect 3234 3168 3238 3172
rect 3252 3168 3256 3172
rect 3274 3165 3278 3169
rect 3299 3165 3303 3169
rect 3309 3168 3313 3172
rect 3325 3168 3329 3172
rect 3345 3165 3349 3169
rect 3352 3168 3356 3172
rect 3145 3158 3149 3162
rect 3184 3158 3188 3162
rect 3228 3158 3232 3162
rect 3259 3158 3263 3162
rect 3281 3158 3285 3162
rect 3346 3158 3350 3162
rect 1507 3150 1511 3154
rect 1895 3150 1899 3154
rect 1904 3151 1910 3155
rect 1995 3151 1999 3155
rect 2029 3151 2033 3155
rect 2046 3151 2050 3155
rect 2102 3151 2106 3155
rect 2119 3151 2123 3155
rect 2147 3151 2151 3155
rect 2230 3151 2234 3155
rect 2256 3151 2260 3155
rect 2290 3151 2294 3155
rect 2307 3151 2311 3155
rect 2363 3151 2367 3155
rect 2380 3151 2384 3155
rect 2408 3151 2412 3155
rect 2452 3150 2456 3154
rect 2840 3150 2844 3154
rect 2849 3151 2855 3155
rect 2940 3151 2944 3155
rect 2974 3151 2978 3155
rect 2991 3151 2995 3155
rect 3047 3151 3051 3155
rect 3064 3151 3068 3155
rect 3092 3151 3096 3155
rect 3175 3151 3179 3155
rect 3201 3151 3205 3155
rect 3235 3151 3239 3155
rect 3252 3151 3256 3155
rect 3308 3151 3312 3155
rect 3325 3151 3329 3155
rect 3353 3151 3357 3155
rect 1630 3143 1635 3147
rect 1763 3143 1767 3147
rect 1940 3144 1946 3148
rect 2004 3144 2008 3148
rect 2238 3144 2242 3148
rect 2424 3145 2428 3149
rect 2436 3145 2440 3149
rect 2575 3143 2580 3147
rect 2708 3143 2712 3147
rect 2885 3144 2891 3148
rect 2949 3144 2953 3148
rect 3183 3144 3187 3148
rect 3369 3145 3373 3149
rect 3381 3145 3385 3149
rect 1638 3136 1642 3140
rect 1928 3136 1934 3140
rect 2248 3137 2252 3141
rect 2413 3137 2417 3141
rect 1622 3131 1626 3135
rect 1654 3131 1658 3135
rect 1976 3130 1982 3134
rect 2583 3136 2587 3140
rect 2873 3136 2879 3140
rect 3193 3137 3197 3141
rect 3358 3137 3362 3141
rect 2567 3131 2571 3135
rect 2599 3131 2603 3135
rect 2921 3130 2927 3134
rect 1491 3123 1495 3127
rect 1622 3123 1626 3127
rect 1654 3123 1658 3127
rect 2567 3123 2571 3127
rect 2599 3123 2603 3127
rect 1638 3116 1642 3120
rect 1895 3116 1899 3120
rect 1964 3116 1970 3120
rect 2296 3116 2300 3120
rect 2332 3116 2336 3120
rect 2399 3116 2403 3120
rect 2583 3116 2587 3120
rect 2840 3116 2844 3120
rect 2909 3116 2915 3120
rect 3241 3116 3245 3120
rect 3277 3116 3281 3120
rect 3344 3116 3348 3120
rect 1895 3108 1899 3112
rect 1904 3109 1910 3113
rect 2282 3109 2286 3113
rect 1622 3104 1626 3108
rect 1654 3104 1658 3108
rect 1638 3100 1642 3104
rect 2296 3102 2300 3106
rect 2346 3102 2350 3106
rect 2399 3102 2403 3106
rect 2840 3108 2844 3112
rect 2849 3109 2855 3113
rect 3227 3109 3231 3113
rect 2567 3104 2571 3108
rect 2599 3104 2603 3108
rect 2583 3100 2587 3104
rect 3241 3102 3245 3106
rect 3291 3102 3295 3106
rect 3344 3102 3348 3106
rect 1630 3093 1635 3097
rect 1764 3093 1768 3097
rect 2319 3091 2323 3095
rect 1513 3086 1517 3090
rect 1549 3086 1553 3090
rect 1616 3086 1620 3090
rect 1645 3086 1649 3090
rect 1681 3086 1685 3090
rect 1748 3086 1752 3090
rect 1777 3086 1781 3090
rect 1813 3086 1817 3090
rect 1880 3086 1884 3090
rect 1964 3086 1970 3090
rect 1904 3079 1910 3083
rect 2290 3082 2294 3086
rect 2303 3085 2307 3091
rect 2340 3085 2344 3091
rect 2353 3087 2357 3091
rect 2377 3091 2381 3095
rect 2575 3093 2580 3097
rect 2709 3093 2713 3097
rect 3264 3091 3268 3095
rect 2361 3085 2365 3091
rect 2398 3085 2402 3091
rect 2414 3085 2418 3091
rect 2458 3086 2462 3090
rect 2494 3086 2498 3090
rect 2561 3086 2565 3090
rect 2590 3086 2594 3090
rect 2626 3086 2630 3090
rect 2693 3086 2697 3090
rect 2722 3086 2726 3090
rect 2758 3086 2762 3090
rect 2825 3086 2829 3090
rect 2909 3086 2915 3090
rect 1513 3072 1517 3076
rect 1563 3072 1567 3076
rect 1616 3072 1620 3076
rect 1645 3072 1649 3076
rect 1695 3072 1699 3076
rect 1748 3072 1752 3076
rect 1777 3072 1781 3076
rect 1827 3072 1831 3076
rect 1880 3072 1884 3076
rect 2303 3072 2307 3076
rect 2319 3072 2323 3078
rect 2353 3078 2357 3082
rect 2340 3072 2344 3076
rect 1536 3061 1540 3065
rect 1507 3052 1511 3056
rect 1520 3055 1524 3061
rect 1557 3055 1561 3061
rect 1570 3057 1574 3061
rect 1594 3061 1598 3065
rect 1668 3061 1672 3065
rect 1578 3055 1582 3061
rect 1615 3055 1619 3061
rect 1631 3055 1635 3061
rect 1652 3055 1656 3061
rect 1689 3055 1693 3061
rect 1702 3057 1706 3061
rect 1726 3061 1730 3065
rect 1800 3061 1804 3065
rect 1710 3055 1714 3061
rect 1747 3055 1751 3061
rect 1763 3055 1767 3061
rect 1784 3055 1788 3061
rect 1821 3055 1825 3061
rect 1834 3057 1838 3061
rect 1858 3061 1862 3065
rect 1842 3055 1846 3061
rect 1879 3055 1883 3061
rect 1895 3057 1899 3061
rect 2361 3072 2365 3076
rect 2377 3072 2381 3078
rect 2849 3079 2855 3083
rect 3235 3082 3239 3086
rect 3248 3085 3252 3091
rect 3285 3085 3289 3091
rect 3298 3087 3302 3091
rect 3322 3091 3326 3095
rect 3306 3085 3310 3091
rect 3343 3085 3347 3091
rect 3359 3085 3363 3091
rect 2398 3072 2402 3076
rect 2414 3072 2418 3076
rect 2458 3072 2462 3076
rect 2508 3072 2512 3076
rect 2561 3072 2565 3076
rect 2590 3072 2594 3076
rect 2640 3072 2644 3076
rect 2693 3072 2697 3076
rect 2722 3072 2726 3076
rect 2772 3072 2776 3076
rect 2825 3072 2829 3076
rect 3248 3072 3252 3076
rect 3264 3072 3268 3078
rect 3298 3078 3302 3082
rect 3285 3072 3289 3076
rect 2296 3061 2300 3065
rect 2333 3059 2337 3063
rect 2353 3059 2357 3063
rect 2397 3059 2401 3063
rect 2481 3061 2485 3065
rect 1520 3042 1524 3046
rect 1536 3042 1540 3048
rect 1570 3048 1574 3052
rect 1557 3042 1561 3046
rect 1578 3042 1582 3046
rect 1594 3042 1598 3048
rect 1615 3042 1619 3046
rect 1631 3042 1635 3046
rect 1652 3042 1656 3046
rect 1668 3042 1672 3048
rect 1702 3048 1706 3052
rect 1689 3042 1693 3046
rect 1710 3042 1714 3046
rect 1726 3042 1730 3048
rect 1747 3042 1751 3046
rect 1763 3042 1767 3046
rect 1784 3042 1788 3046
rect 1800 3042 1804 3048
rect 1834 3048 1838 3052
rect 1821 3042 1825 3046
rect 1842 3042 1846 3046
rect 1858 3042 1862 3048
rect 1916 3052 1922 3056
rect 2452 3052 2456 3056
rect 2465 3055 2469 3061
rect 2502 3055 2506 3061
rect 2515 3057 2519 3061
rect 2539 3061 2543 3065
rect 2613 3061 2617 3065
rect 2523 3055 2527 3061
rect 2560 3055 2564 3061
rect 2576 3055 2580 3061
rect 2597 3055 2601 3061
rect 2634 3055 2638 3061
rect 2647 3057 2651 3061
rect 2671 3061 2675 3065
rect 2745 3061 2749 3065
rect 2655 3055 2659 3061
rect 2692 3055 2696 3061
rect 2708 3055 2712 3061
rect 2729 3055 2733 3061
rect 2766 3055 2770 3061
rect 2779 3057 2783 3061
rect 2803 3061 2807 3065
rect 2787 3055 2791 3061
rect 2824 3055 2828 3061
rect 2840 3057 2844 3061
rect 3306 3072 3310 3076
rect 3322 3072 3326 3078
rect 3343 3072 3347 3076
rect 3359 3072 3363 3076
rect 3241 3061 3245 3065
rect 3278 3059 3282 3063
rect 3298 3059 3302 3063
rect 3342 3059 3346 3063
rect 1879 3042 1883 3046
rect 1895 3042 1899 3046
rect 1952 3045 1958 3049
rect 2296 3045 2300 3049
rect 2347 3045 2351 3049
rect 2397 3045 2401 3049
rect 2465 3042 2469 3046
rect 2481 3042 2485 3048
rect 2515 3048 2519 3052
rect 2502 3042 2506 3046
rect 1513 3031 1517 3035
rect 1550 3029 1554 3033
rect 1570 3029 1574 3033
rect 1614 3029 1618 3033
rect 1645 3031 1649 3035
rect 1682 3029 1686 3033
rect 1702 3029 1706 3033
rect 1746 3029 1750 3033
rect 1777 3031 1781 3035
rect 1814 3029 1818 3033
rect 1834 3029 1838 3033
rect 1878 3029 1882 3033
rect 2289 3037 2293 3041
rect 2414 3038 2418 3042
rect 2523 3042 2527 3046
rect 2539 3042 2543 3048
rect 2560 3042 2564 3046
rect 2576 3042 2580 3046
rect 2597 3042 2601 3046
rect 2613 3042 2617 3048
rect 2647 3048 2651 3052
rect 2634 3042 2638 3046
rect 2655 3042 2659 3046
rect 2671 3042 2675 3048
rect 2692 3042 2696 3046
rect 2708 3042 2712 3046
rect 2729 3042 2733 3046
rect 2745 3042 2749 3048
rect 2779 3048 2783 3052
rect 2766 3042 2770 3046
rect 2787 3042 2791 3046
rect 2803 3042 2807 3048
rect 2861 3052 2867 3056
rect 2824 3042 2828 3046
rect 2840 3042 2844 3046
rect 2897 3045 2903 3049
rect 3241 3045 3245 3049
rect 3292 3045 3296 3049
rect 3342 3045 3346 3049
rect 1964 3030 1970 3034
rect 2296 3030 2300 3034
rect 2332 3030 2336 3034
rect 2399 3030 2403 3034
rect 1916 3022 1922 3026
rect 2282 3023 2286 3027
rect 2458 3031 2462 3035
rect 2495 3029 2499 3033
rect 2515 3029 2519 3033
rect 2559 3029 2563 3033
rect 2590 3031 2594 3035
rect 2627 3029 2631 3033
rect 2647 3029 2651 3033
rect 2691 3029 2695 3033
rect 2722 3031 2726 3035
rect 2759 3029 2763 3033
rect 2779 3029 2783 3033
rect 2823 3029 2827 3033
rect 3234 3037 3238 3041
rect 3359 3038 3363 3042
rect 2909 3030 2915 3034
rect 3241 3030 3245 3034
rect 3277 3030 3281 3034
rect 3344 3030 3348 3034
rect 1513 3015 1517 3019
rect 1564 3015 1568 3019
rect 1614 3015 1618 3019
rect 1645 3015 1649 3019
rect 1696 3015 1700 3019
rect 1746 3015 1750 3019
rect 1777 3015 1781 3019
rect 1828 3015 1832 3019
rect 1878 3015 1882 3019
rect 1952 3015 1958 3019
rect 2296 3016 2300 3020
rect 2346 3016 2350 3020
rect 2399 3016 2403 3020
rect 2861 3022 2867 3026
rect 3227 3023 3231 3027
rect 2458 3015 2462 3019
rect 2509 3015 2513 3019
rect 2559 3015 2563 3019
rect 2590 3015 2594 3019
rect 2641 3015 2645 3019
rect 2691 3015 2695 3019
rect 2722 3015 2726 3019
rect 2773 3015 2777 3019
rect 2823 3015 2827 3019
rect 2897 3015 2903 3019
rect 3241 3016 3245 3020
rect 3291 3016 3295 3020
rect 3344 3016 3348 3020
rect 1506 3008 1510 3012
rect 1895 3008 1899 3012
rect 2319 3005 2323 3009
rect 1513 3000 1517 3004
rect 1549 3000 1553 3004
rect 1616 3000 1620 3004
rect 1645 3000 1649 3004
rect 1681 3000 1685 3004
rect 1748 3000 1752 3004
rect 1777 3000 1781 3004
rect 1813 3000 1817 3004
rect 1880 3000 1884 3004
rect 1964 3000 1970 3004
rect 1904 2993 1910 2997
rect 2290 2996 2294 3000
rect 2303 2999 2307 3005
rect 2340 2999 2344 3005
rect 2353 3001 2357 3005
rect 2377 3005 2381 3009
rect 2451 3008 2455 3012
rect 2840 3008 2844 3012
rect 3264 3005 3268 3009
rect 2361 2999 2365 3005
rect 2398 2999 2402 3005
rect 2414 3001 2418 3005
rect 2436 2999 2440 3003
rect 2458 3000 2462 3004
rect 2494 3000 2498 3004
rect 2561 3000 2565 3004
rect 2590 3000 2594 3004
rect 2626 3000 2630 3004
rect 2693 3000 2697 3004
rect 2722 3000 2726 3004
rect 2758 3000 2762 3004
rect 2825 3000 2829 3004
rect 2909 3000 2915 3004
rect 1513 2986 1517 2990
rect 1563 2986 1567 2990
rect 1616 2986 1620 2990
rect 1645 2986 1649 2990
rect 1695 2986 1699 2990
rect 1748 2986 1752 2990
rect 1777 2986 1781 2990
rect 1827 2986 1831 2990
rect 1880 2986 1884 2990
rect 2303 2986 2307 2990
rect 2319 2986 2323 2992
rect 2353 2992 2357 2996
rect 2340 2986 2344 2990
rect 1536 2975 1540 2979
rect 1507 2966 1511 2970
rect 1520 2969 1524 2975
rect 1557 2969 1561 2975
rect 1570 2971 1574 2975
rect 1594 2975 1598 2979
rect 1668 2975 1672 2979
rect 1578 2969 1582 2975
rect 1615 2969 1619 2975
rect 1631 2969 1635 2975
rect 1652 2969 1656 2975
rect 1689 2969 1693 2975
rect 1702 2971 1706 2975
rect 1726 2975 1730 2979
rect 1800 2975 1804 2979
rect 1710 2969 1714 2975
rect 1747 2969 1751 2975
rect 1763 2969 1767 2975
rect 1784 2969 1788 2975
rect 1821 2969 1825 2975
rect 1834 2971 1838 2975
rect 1858 2975 1862 2979
rect 1842 2969 1846 2975
rect 1879 2969 1883 2975
rect 1895 2971 1899 2975
rect 2361 2986 2365 2990
rect 2377 2986 2381 2992
rect 2398 2986 2402 2990
rect 2414 2986 2418 2995
rect 2849 2993 2855 2997
rect 3235 2996 3239 3000
rect 3248 2999 3252 3005
rect 3285 2999 3289 3005
rect 3298 3001 3302 3005
rect 3322 3005 3326 3009
rect 3306 2999 3310 3005
rect 3343 2999 3347 3005
rect 3359 3001 3363 3005
rect 3381 2999 3385 3003
rect 2436 2983 2440 2987
rect 2458 2986 2462 2990
rect 2508 2986 2512 2990
rect 2561 2986 2565 2990
rect 2590 2986 2594 2990
rect 2640 2986 2644 2990
rect 2693 2986 2697 2990
rect 2722 2986 2726 2990
rect 2772 2986 2776 2990
rect 2825 2986 2829 2990
rect 3248 2986 3252 2990
rect 3264 2986 3268 2992
rect 3298 2992 3302 2996
rect 3285 2986 3289 2990
rect 2296 2975 2300 2979
rect 2333 2973 2337 2977
rect 2353 2973 2357 2977
rect 2397 2973 2401 2977
rect 2481 2975 2485 2979
rect 1520 2956 1524 2960
rect 1536 2956 1540 2962
rect 1570 2962 1574 2966
rect 1557 2956 1561 2960
rect 1578 2956 1582 2960
rect 1594 2956 1598 2962
rect 1615 2956 1619 2960
rect 1631 2956 1635 2960
rect 1652 2956 1656 2960
rect 1668 2956 1672 2962
rect 1702 2962 1706 2966
rect 1689 2956 1693 2960
rect 1710 2956 1714 2960
rect 1726 2956 1730 2962
rect 1747 2956 1751 2960
rect 1763 2956 1767 2960
rect 1784 2956 1788 2960
rect 1800 2956 1804 2962
rect 1834 2962 1838 2966
rect 1821 2956 1825 2960
rect 1842 2956 1846 2960
rect 1858 2956 1862 2962
rect 1916 2966 1922 2970
rect 2452 2966 2456 2970
rect 2465 2969 2469 2975
rect 2502 2969 2506 2975
rect 2515 2971 2519 2975
rect 2539 2975 2543 2979
rect 2613 2975 2617 2979
rect 2523 2969 2527 2975
rect 2560 2969 2564 2975
rect 2576 2969 2580 2975
rect 2597 2969 2601 2975
rect 2634 2969 2638 2975
rect 2647 2971 2651 2975
rect 2671 2975 2675 2979
rect 2745 2975 2749 2979
rect 2655 2969 2659 2975
rect 2692 2969 2696 2975
rect 2708 2969 2712 2975
rect 2729 2969 2733 2975
rect 2766 2969 2770 2975
rect 2779 2971 2783 2975
rect 2803 2975 2807 2979
rect 2787 2969 2791 2975
rect 2824 2969 2828 2975
rect 2840 2971 2844 2975
rect 3306 2986 3310 2990
rect 3322 2986 3326 2992
rect 3343 2986 3347 2990
rect 3359 2986 3363 2995
rect 3381 2983 3385 2987
rect 3241 2975 3245 2979
rect 3278 2973 3282 2977
rect 3298 2973 3302 2977
rect 3342 2973 3346 2977
rect 1879 2956 1883 2960
rect 1895 2956 1899 2960
rect 1952 2959 1958 2963
rect 2296 2959 2300 2963
rect 2347 2959 2351 2963
rect 2397 2959 2401 2963
rect 2465 2956 2469 2960
rect 2481 2956 2485 2962
rect 2515 2962 2519 2966
rect 2502 2956 2506 2960
rect 2523 2956 2527 2960
rect 2539 2956 2543 2962
rect 2560 2956 2564 2960
rect 2576 2956 2580 2960
rect 2597 2956 2601 2960
rect 2613 2956 2617 2962
rect 2647 2962 2651 2966
rect 2634 2956 2638 2960
rect 2655 2956 2659 2960
rect 2671 2956 2675 2962
rect 2692 2956 2696 2960
rect 2708 2956 2712 2960
rect 2729 2956 2733 2960
rect 2745 2956 2749 2962
rect 2779 2962 2783 2966
rect 2766 2956 2770 2960
rect 2787 2956 2791 2960
rect 2803 2956 2807 2962
rect 2861 2966 2867 2970
rect 2824 2956 2828 2960
rect 2840 2956 2844 2960
rect 2897 2959 2903 2963
rect 3241 2959 3245 2963
rect 3292 2959 3296 2963
rect 3342 2959 3346 2963
rect 1513 2945 1517 2949
rect 1550 2943 1554 2947
rect 1570 2943 1574 2947
rect 1614 2943 1618 2947
rect 1645 2945 1649 2949
rect 1682 2943 1686 2947
rect 1702 2943 1706 2947
rect 1746 2943 1750 2947
rect 1777 2945 1781 2949
rect 1814 2943 1818 2947
rect 1834 2943 1838 2947
rect 1878 2943 1882 2947
rect 2458 2945 2462 2949
rect 2495 2943 2499 2947
rect 2515 2943 2519 2947
rect 2559 2943 2563 2947
rect 2590 2945 2594 2949
rect 2627 2943 2631 2947
rect 2647 2943 2651 2947
rect 2691 2943 2695 2947
rect 2722 2945 2726 2949
rect 2759 2943 2763 2947
rect 2779 2943 2783 2947
rect 2823 2943 2827 2947
rect 1916 2936 1922 2940
rect 2861 2936 2867 2940
rect 1513 2929 1517 2933
rect 1564 2929 1568 2933
rect 1614 2929 1618 2933
rect 1645 2929 1649 2933
rect 1696 2929 1700 2933
rect 1746 2929 1750 2933
rect 1777 2929 1781 2933
rect 1828 2929 1832 2933
rect 1878 2929 1882 2933
rect 1952 2929 1958 2933
rect 2458 2929 2462 2933
rect 2509 2929 2513 2933
rect 2559 2929 2563 2933
rect 2590 2929 2594 2933
rect 2641 2929 2645 2933
rect 2691 2929 2695 2933
rect 2722 2929 2726 2933
rect 2773 2929 2777 2933
rect 2823 2929 2827 2933
rect 2897 2929 2903 2933
rect 1506 2922 1510 2926
rect 1895 2922 1899 2926
rect 2451 2922 2455 2926
rect 2840 2922 2844 2926
rect 1631 2915 1635 2919
rect 1739 2915 1743 2919
rect 1763 2915 1767 2919
rect 2576 2915 2580 2919
rect 2684 2915 2688 2919
rect 2708 2915 2712 2919
rect 1755 2908 1759 2912
rect 1739 2904 1743 2908
rect 1771 2904 1775 2908
rect 2700 2908 2704 2912
rect 2684 2904 2688 2908
rect 2716 2904 2720 2908
rect 1739 2897 1743 2901
rect 1771 2897 1775 2901
rect 2436 2897 2440 2901
rect 2684 2897 2688 2901
rect 2716 2897 2720 2901
rect 3381 2897 3385 2901
rect 1755 2890 1759 2894
rect 1895 2890 1899 2894
rect 2700 2890 2704 2894
rect 2840 2890 2844 2894
rect 1895 2882 1899 2886
rect 2840 2882 2844 2886
rect 1739 2878 1743 2882
rect 1771 2878 1775 2882
rect 1755 2874 1759 2878
rect 2684 2878 2688 2882
rect 2716 2878 2720 2882
rect 2700 2874 2704 2878
rect 1631 2867 1635 2871
rect 1739 2867 1743 2871
rect 1763 2867 1767 2871
rect 2576 2867 2580 2871
rect 2684 2867 2688 2871
rect 2708 2867 2712 2871
rect 1513 2860 1517 2864
rect 1549 2860 1553 2864
rect 1616 2860 1620 2864
rect 1645 2860 1649 2864
rect 1681 2860 1685 2864
rect 1748 2860 1752 2864
rect 1777 2860 1781 2864
rect 1813 2860 1817 2864
rect 1880 2860 1884 2864
rect 1964 2860 1970 2864
rect 2458 2860 2462 2864
rect 2494 2860 2498 2864
rect 2561 2860 2565 2864
rect 2590 2860 2594 2864
rect 2626 2860 2630 2864
rect 2693 2860 2697 2864
rect 2722 2860 2726 2864
rect 2758 2860 2762 2864
rect 2825 2860 2829 2864
rect 2909 2860 2915 2864
rect 1904 2853 1910 2857
rect 2849 2853 2855 2857
rect 1513 2846 1517 2850
rect 1563 2846 1567 2850
rect 1616 2846 1620 2850
rect 1645 2846 1649 2850
rect 1695 2846 1699 2850
rect 1748 2846 1752 2850
rect 1777 2846 1781 2850
rect 1827 2846 1831 2850
rect 1880 2846 1884 2850
rect 2458 2846 2462 2850
rect 2508 2846 2512 2850
rect 2561 2846 2565 2850
rect 2590 2846 2594 2850
rect 2640 2846 2644 2850
rect 2693 2846 2697 2850
rect 2722 2846 2726 2850
rect 2772 2846 2776 2850
rect 2825 2846 2829 2850
rect 1536 2835 1540 2839
rect 1507 2826 1511 2830
rect 1520 2829 1524 2835
rect 1557 2829 1561 2835
rect 1570 2831 1574 2835
rect 1594 2835 1598 2839
rect 1668 2835 1672 2839
rect 1578 2829 1582 2835
rect 1615 2829 1619 2835
rect 1631 2829 1635 2835
rect 1652 2829 1656 2835
rect 1689 2829 1693 2835
rect 1702 2831 1706 2835
rect 1726 2835 1730 2839
rect 1800 2835 1804 2839
rect 1710 2829 1714 2835
rect 1747 2829 1751 2835
rect 1763 2829 1767 2835
rect 1784 2829 1788 2835
rect 1821 2829 1825 2835
rect 1834 2831 1838 2835
rect 1858 2835 1862 2839
rect 2481 2835 2485 2839
rect 1842 2829 1846 2835
rect 1879 2829 1883 2835
rect 1895 2831 1899 2835
rect 1520 2816 1524 2820
rect 1536 2816 1540 2822
rect 1570 2822 1574 2826
rect 1557 2816 1561 2820
rect 1578 2816 1582 2820
rect 1594 2816 1598 2822
rect 1615 2816 1619 2820
rect 1631 2816 1635 2820
rect 1652 2816 1656 2820
rect 1668 2816 1672 2822
rect 1702 2822 1706 2826
rect 1689 2816 1693 2820
rect 1710 2816 1714 2820
rect 1726 2816 1730 2822
rect 1747 2816 1751 2820
rect 1763 2816 1767 2820
rect 1784 2816 1788 2820
rect 1800 2816 1804 2822
rect 1834 2822 1838 2826
rect 1821 2816 1825 2820
rect 1842 2816 1846 2820
rect 1858 2816 1862 2822
rect 2452 2826 2456 2830
rect 2465 2829 2469 2835
rect 2502 2829 2506 2835
rect 2515 2831 2519 2835
rect 2539 2835 2543 2839
rect 2613 2835 2617 2839
rect 2523 2829 2527 2835
rect 2560 2829 2564 2835
rect 2576 2829 2580 2835
rect 2597 2829 2601 2835
rect 2634 2829 2638 2835
rect 2647 2831 2651 2835
rect 2671 2835 2675 2839
rect 2745 2835 2749 2839
rect 2655 2829 2659 2835
rect 2692 2829 2696 2835
rect 2708 2829 2712 2835
rect 2729 2829 2733 2835
rect 2766 2829 2770 2835
rect 2779 2831 2783 2835
rect 2803 2835 2807 2839
rect 2787 2829 2791 2835
rect 2824 2829 2828 2835
rect 2840 2831 2844 2835
rect 1879 2816 1883 2820
rect 1895 2816 1899 2820
rect 2465 2816 2469 2820
rect 2481 2816 2485 2822
rect 2515 2822 2519 2826
rect 2502 2816 2506 2820
rect 2523 2816 2527 2820
rect 2539 2816 2543 2822
rect 2560 2816 2564 2820
rect 2576 2816 2580 2820
rect 2597 2816 2601 2820
rect 2613 2816 2617 2822
rect 2647 2822 2651 2826
rect 2634 2816 2638 2820
rect 2655 2816 2659 2820
rect 2671 2816 2675 2822
rect 2692 2816 2696 2820
rect 2708 2816 2712 2820
rect 2729 2816 2733 2820
rect 2745 2816 2749 2822
rect 2779 2822 2783 2826
rect 2766 2816 2770 2820
rect 2787 2816 2791 2820
rect 2803 2816 2807 2822
rect 2824 2816 2828 2820
rect 2840 2816 2844 2820
rect 1513 2805 1517 2809
rect 1550 2803 1554 2807
rect 1570 2803 1574 2807
rect 1614 2803 1618 2807
rect 1645 2805 1649 2809
rect 1682 2803 1686 2807
rect 1702 2803 1706 2807
rect 1746 2803 1750 2807
rect 1777 2805 1781 2809
rect 1814 2803 1818 2807
rect 1834 2803 1838 2807
rect 1878 2803 1882 2807
rect 2458 2805 2462 2809
rect 2495 2803 2499 2807
rect 2515 2803 2519 2807
rect 2559 2803 2563 2807
rect 2590 2805 2594 2809
rect 2627 2803 2631 2807
rect 2647 2803 2651 2807
rect 2691 2803 2695 2807
rect 2722 2805 2726 2809
rect 2759 2803 2763 2807
rect 2779 2803 2783 2807
rect 2823 2803 2827 2807
rect 1916 2796 1922 2800
rect 2861 2796 2867 2800
rect 1513 2789 1517 2793
rect 1564 2789 1568 2793
rect 1614 2789 1618 2793
rect 1645 2789 1649 2793
rect 1696 2789 1700 2793
rect 1746 2789 1750 2793
rect 1777 2789 1781 2793
rect 1828 2789 1832 2793
rect 1878 2789 1882 2793
rect 1952 2789 1958 2793
rect 2458 2789 2462 2793
rect 2509 2789 2513 2793
rect 2559 2789 2563 2793
rect 2590 2789 2594 2793
rect 2641 2789 2645 2793
rect 2691 2789 2695 2793
rect 2722 2789 2726 2793
rect 2773 2789 2777 2793
rect 2823 2789 2827 2793
rect 2897 2789 2903 2793
rect 1964 2781 1970 2785
rect 1997 2781 2001 2785
rect 2033 2781 2037 2785
rect 2100 2781 2104 2785
rect 2129 2781 2133 2785
rect 2165 2781 2169 2785
rect 2232 2781 2236 2785
rect 2261 2781 2265 2785
rect 2297 2781 2301 2785
rect 2364 2781 2368 2785
rect 2393 2781 2397 2785
rect 2429 2781 2433 2785
rect 2496 2781 2500 2785
rect 2909 2781 2915 2785
rect 2942 2781 2946 2785
rect 2978 2781 2982 2785
rect 3045 2781 3049 2785
rect 3074 2781 3078 2785
rect 3110 2781 3114 2785
rect 3177 2781 3181 2785
rect 3206 2781 3210 2785
rect 3242 2781 3246 2785
rect 3309 2781 3313 2785
rect 3338 2781 3342 2785
rect 3374 2781 3378 2785
rect 3441 2781 3445 2785
rect 1904 2774 1910 2778
rect 2849 2774 2855 2778
rect 1997 2767 2001 2771
rect 2047 2767 2051 2771
rect 2100 2767 2104 2771
rect 2129 2767 2133 2771
rect 2179 2767 2183 2771
rect 2232 2767 2236 2771
rect 2261 2767 2265 2771
rect 2311 2767 2315 2771
rect 2364 2767 2368 2771
rect 2393 2767 2397 2771
rect 2443 2767 2447 2771
rect 2496 2767 2500 2771
rect 2942 2767 2946 2771
rect 2992 2767 2996 2771
rect 3045 2767 3049 2771
rect 3074 2767 3078 2771
rect 3124 2767 3128 2771
rect 3177 2767 3181 2771
rect 3206 2767 3210 2771
rect 3256 2767 3260 2771
rect 3309 2767 3313 2771
rect 3338 2767 3342 2771
rect 3388 2767 3392 2771
rect 3441 2767 3445 2771
rect 2020 2756 2024 2760
rect 1645 2748 1649 2752
rect 1681 2748 1685 2752
rect 1748 2748 1752 2752
rect 1964 2748 1970 2752
rect 1991 2747 1995 2751
rect 2004 2750 2008 2756
rect 2041 2750 2045 2756
rect 2054 2752 2058 2756
rect 2078 2756 2082 2760
rect 2152 2756 2156 2760
rect 2062 2750 2066 2756
rect 2099 2750 2103 2756
rect 2115 2752 2119 2756
rect 1904 2741 1910 2745
rect 1645 2734 1649 2738
rect 1695 2734 1699 2738
rect 1748 2734 1752 2738
rect 2004 2737 2008 2741
rect 2020 2737 2024 2743
rect 2054 2743 2058 2747
rect 2041 2737 2045 2741
rect 2062 2737 2066 2741
rect 2078 2737 2082 2743
rect 2123 2747 2127 2751
rect 2136 2750 2140 2756
rect 2173 2750 2177 2756
rect 2186 2752 2190 2756
rect 2210 2756 2214 2760
rect 2284 2756 2288 2760
rect 2194 2750 2198 2756
rect 2231 2750 2235 2756
rect 2247 2752 2251 2756
rect 2099 2737 2103 2741
rect 2115 2737 2119 2741
rect 2136 2737 2140 2741
rect 2152 2737 2156 2743
rect 2186 2743 2190 2747
rect 2173 2737 2177 2741
rect 2194 2737 2198 2741
rect 2210 2737 2214 2743
rect 2255 2747 2259 2751
rect 2268 2750 2272 2756
rect 2305 2750 2309 2756
rect 2318 2752 2322 2756
rect 2342 2756 2346 2760
rect 2416 2756 2420 2760
rect 2326 2750 2330 2756
rect 2363 2750 2367 2756
rect 2379 2752 2383 2756
rect 2231 2737 2235 2741
rect 2247 2737 2251 2741
rect 2268 2737 2272 2741
rect 2284 2737 2288 2743
rect 2318 2743 2322 2747
rect 2305 2737 2309 2741
rect 2326 2737 2330 2741
rect 2342 2737 2346 2743
rect 2387 2747 2391 2751
rect 2400 2750 2404 2756
rect 2437 2750 2441 2756
rect 2450 2752 2454 2756
rect 2474 2756 2478 2760
rect 2965 2756 2969 2760
rect 2458 2750 2462 2756
rect 2495 2750 2499 2756
rect 2511 2752 2515 2756
rect 2590 2748 2594 2752
rect 2626 2748 2630 2752
rect 2693 2748 2697 2752
rect 2909 2748 2915 2752
rect 2363 2737 2367 2741
rect 2379 2737 2383 2741
rect 2400 2737 2404 2741
rect 2416 2737 2420 2743
rect 2450 2743 2454 2747
rect 2437 2737 2441 2741
rect 1668 2723 1672 2727
rect 1630 2714 1634 2718
rect 1652 2717 1656 2723
rect 1689 2717 1693 2723
rect 1702 2719 1706 2723
rect 1726 2723 1730 2727
rect 1710 2717 1714 2723
rect 1747 2717 1751 2723
rect 1763 2717 1767 2723
rect 1997 2726 2001 2730
rect 2034 2724 2038 2728
rect 2054 2724 2058 2728
rect 2098 2724 2102 2728
rect 2129 2726 2133 2730
rect 2166 2724 2170 2728
rect 2186 2724 2190 2728
rect 2230 2724 2234 2728
rect 2261 2726 2265 2730
rect 2298 2724 2302 2728
rect 2318 2724 2322 2728
rect 2362 2724 2366 2728
rect 2379 2729 2383 2733
rect 2458 2737 2462 2741
rect 2474 2737 2478 2743
rect 2936 2747 2940 2751
rect 2949 2750 2953 2756
rect 2986 2750 2990 2756
rect 2999 2752 3003 2756
rect 3023 2756 3027 2760
rect 3097 2756 3101 2760
rect 3007 2750 3011 2756
rect 3044 2750 3048 2756
rect 3060 2752 3064 2756
rect 2849 2741 2855 2745
rect 2495 2737 2499 2741
rect 2511 2737 2515 2741
rect 2393 2726 2397 2730
rect 2430 2724 2434 2728
rect 2450 2724 2454 2728
rect 2494 2724 2498 2728
rect 2511 2729 2515 2733
rect 2590 2734 2594 2738
rect 2640 2734 2644 2738
rect 2693 2734 2697 2738
rect 2949 2737 2953 2741
rect 2965 2737 2969 2743
rect 2999 2743 3003 2747
rect 2986 2737 2990 2741
rect 3007 2737 3011 2741
rect 3023 2737 3027 2743
rect 3068 2747 3072 2751
rect 3081 2750 3085 2756
rect 3118 2750 3122 2756
rect 3131 2752 3135 2756
rect 3155 2756 3159 2760
rect 3229 2756 3233 2760
rect 3139 2750 3143 2756
rect 3176 2750 3180 2756
rect 3192 2752 3196 2756
rect 3044 2737 3048 2741
rect 3060 2737 3064 2741
rect 3081 2737 3085 2741
rect 3097 2737 3101 2743
rect 3131 2743 3135 2747
rect 3118 2737 3122 2741
rect 3139 2737 3143 2741
rect 3155 2737 3159 2743
rect 3200 2747 3204 2751
rect 3213 2750 3217 2756
rect 3250 2750 3254 2756
rect 3263 2752 3267 2756
rect 3287 2756 3291 2760
rect 3361 2756 3365 2760
rect 3271 2750 3275 2756
rect 3308 2750 3312 2756
rect 3324 2752 3328 2756
rect 3176 2737 3180 2741
rect 3192 2737 3196 2741
rect 3213 2737 3217 2741
rect 3229 2737 3233 2743
rect 3263 2743 3267 2747
rect 3250 2737 3254 2741
rect 3271 2737 3275 2741
rect 3287 2737 3291 2743
rect 3332 2747 3336 2751
rect 3345 2750 3349 2756
rect 3382 2750 3386 2756
rect 3395 2752 3399 2756
rect 3419 2756 3423 2760
rect 3403 2750 3407 2756
rect 3440 2750 3444 2756
rect 3456 2752 3460 2756
rect 3308 2737 3312 2741
rect 3324 2737 3328 2741
rect 3345 2737 3349 2741
rect 3361 2737 3365 2743
rect 3395 2743 3399 2747
rect 3382 2737 3386 2741
rect 2613 2723 2617 2727
rect 1916 2717 1922 2721
rect 1652 2704 1656 2708
rect 1668 2704 1672 2710
rect 1702 2710 1706 2714
rect 1689 2704 1693 2708
rect 1710 2704 1714 2708
rect 1726 2704 1730 2710
rect 2575 2714 2579 2718
rect 2597 2717 2601 2723
rect 2634 2717 2638 2723
rect 2647 2719 2651 2723
rect 2671 2723 2675 2727
rect 2655 2717 2659 2723
rect 2692 2717 2696 2723
rect 2708 2717 2712 2723
rect 2942 2726 2946 2730
rect 2979 2724 2983 2728
rect 2999 2724 3003 2728
rect 3043 2724 3047 2728
rect 3074 2726 3078 2730
rect 3111 2724 3115 2728
rect 3131 2724 3135 2728
rect 3175 2724 3179 2728
rect 3206 2726 3210 2730
rect 3243 2724 3247 2728
rect 3263 2724 3267 2728
rect 3307 2724 3311 2728
rect 3324 2729 3328 2733
rect 3403 2737 3407 2741
rect 3419 2737 3423 2743
rect 3440 2737 3444 2741
rect 3456 2737 3460 2741
rect 3338 2726 3342 2730
rect 3375 2724 3379 2728
rect 3395 2724 3399 2728
rect 3439 2724 3443 2728
rect 3456 2729 3460 2733
rect 2861 2717 2867 2721
rect 1952 2710 1958 2714
rect 1997 2710 2001 2714
rect 2048 2710 2052 2714
rect 2098 2710 2102 2714
rect 2129 2710 2133 2714
rect 2180 2710 2184 2714
rect 2230 2710 2234 2714
rect 2261 2710 2265 2714
rect 2312 2710 2316 2714
rect 2362 2710 2366 2714
rect 2393 2710 2397 2714
rect 2444 2710 2448 2714
rect 2494 2710 2498 2714
rect 1747 2704 1751 2708
rect 1763 2704 1767 2708
rect 2597 2704 2601 2708
rect 2613 2704 2617 2710
rect 2647 2710 2651 2714
rect 2634 2704 2638 2708
rect 1645 2693 1649 2697
rect 1682 2691 1686 2695
rect 1702 2691 1706 2695
rect 1746 2691 1750 2695
rect 1904 2697 1910 2701
rect 1995 2697 1999 2701
rect 2029 2697 2033 2701
rect 2046 2697 2050 2701
rect 2102 2697 2106 2701
rect 2119 2697 2123 2701
rect 2147 2697 2151 2701
rect 2655 2704 2659 2708
rect 2671 2704 2675 2710
rect 2897 2710 2903 2714
rect 2942 2710 2946 2714
rect 2993 2710 2997 2714
rect 3043 2710 3047 2714
rect 3074 2710 3078 2714
rect 3125 2710 3129 2714
rect 3175 2710 3179 2714
rect 3206 2710 3210 2714
rect 3257 2710 3261 2714
rect 3307 2710 3311 2714
rect 3338 2710 3342 2714
rect 3389 2710 3393 2714
rect 3439 2710 3443 2714
rect 2692 2704 2696 2708
rect 2708 2704 2712 2708
rect 1940 2690 1946 2694
rect 2022 2690 2026 2694
rect 2053 2690 2057 2694
rect 2075 2690 2079 2694
rect 2140 2690 2144 2694
rect 1916 2684 1922 2688
rect 1645 2677 1649 2681
rect 1696 2677 1700 2681
rect 1746 2677 1750 2681
rect 1952 2677 1958 2681
rect 1996 2680 2000 2684
rect 2021 2683 2025 2687
rect 2028 2680 2032 2684
rect 2046 2680 2050 2684
rect 2068 2683 2072 2687
rect 2093 2683 2097 2687
rect 2103 2680 2107 2684
rect 2119 2680 2123 2684
rect 2139 2683 2143 2687
rect 2146 2680 2150 2684
rect 2210 2690 2214 2694
rect 1763 2670 1767 2674
rect 1630 2661 1634 2665
rect 1755 2663 1759 2667
rect 1779 2663 1783 2667
rect 1989 2663 1993 2667
rect 1638 2654 1642 2658
rect 1779 2654 1783 2658
rect 2023 2664 2027 2668
rect 2043 2661 2047 2665
rect 2062 2665 2066 2669
rect 2164 2676 2168 2680
rect 2179 2676 2183 2680
rect 2081 2664 2085 2668
rect 2100 2664 2104 2668
rect 2113 2663 2117 2667
rect 2135 2664 2139 2668
rect 2143 2663 2147 2667
rect 2155 2663 2159 2667
rect 1996 2650 2000 2654
rect 2028 2650 2032 2654
rect 2046 2650 2050 2654
rect 2103 2650 2107 2654
rect 2118 2650 2122 2654
rect 2146 2650 2150 2654
rect 1645 2646 1649 2650
rect 1712 2646 1716 2650
rect 1748 2646 1752 2650
rect 1964 2646 1970 2650
rect 2010 2646 2014 2650
rect 2053 2645 2057 2649
rect 2075 2646 2082 2650
rect 2125 2645 2129 2649
rect 1904 2639 1910 2643
rect 1645 2632 1649 2636
rect 1698 2632 1702 2636
rect 1748 2632 1752 2636
rect 1928 2638 1934 2642
rect 2010 2638 2014 2642
rect 2069 2638 2073 2642
rect 2094 2638 2098 2642
rect 2125 2638 2129 2642
rect 2218 2668 2222 2676
rect 2291 2690 2295 2694
rect 2245 2676 2249 2680
rect 2260 2676 2264 2680
rect 2590 2693 2594 2697
rect 2627 2691 2631 2695
rect 2647 2691 2651 2695
rect 2691 2691 2695 2695
rect 2849 2697 2855 2701
rect 2940 2697 2944 2701
rect 2974 2697 2978 2701
rect 2991 2697 2995 2701
rect 3047 2697 3051 2701
rect 3064 2697 3068 2701
rect 3092 2697 3096 2701
rect 2885 2690 2891 2694
rect 2967 2690 2971 2694
rect 2998 2690 3002 2694
rect 3020 2690 3024 2694
rect 3085 2690 3089 2694
rect 2241 2668 2245 2672
rect 2187 2662 2191 2666
rect 2200 2654 2204 2658
rect 2299 2668 2303 2676
rect 2861 2684 2867 2688
rect 2590 2677 2594 2681
rect 2641 2677 2645 2681
rect 2691 2677 2695 2681
rect 2897 2677 2903 2681
rect 2941 2680 2945 2684
rect 2966 2683 2970 2687
rect 2973 2680 2977 2684
rect 2991 2680 2995 2684
rect 3013 2683 3017 2687
rect 3038 2683 3042 2687
rect 3048 2680 3052 2684
rect 3064 2680 3068 2684
rect 3084 2683 3088 2687
rect 3091 2680 3095 2684
rect 3155 2690 3159 2694
rect 2326 2668 2330 2672
rect 2708 2670 2712 2674
rect 2268 2662 2272 2666
rect 2575 2661 2579 2665
rect 2700 2663 2704 2667
rect 2724 2663 2728 2667
rect 2934 2663 2938 2667
rect 2281 2654 2285 2658
rect 2583 2654 2587 2658
rect 2724 2654 2728 2658
rect 2968 2664 2972 2668
rect 2988 2661 2992 2665
rect 3007 2665 3011 2669
rect 3109 2676 3113 2680
rect 3124 2676 3128 2680
rect 3026 2664 3030 2668
rect 3045 2664 3049 2668
rect 3058 2663 3062 2667
rect 3080 2664 3084 2668
rect 3088 2663 3092 2667
rect 3100 2663 3104 2667
rect 2941 2650 2945 2654
rect 2973 2650 2977 2654
rect 2991 2650 2995 2654
rect 3048 2650 3052 2654
rect 3063 2650 3067 2654
rect 3091 2650 3095 2654
rect 2590 2646 2594 2650
rect 2657 2646 2661 2650
rect 2693 2646 2697 2650
rect 2909 2646 2915 2650
rect 2955 2646 2959 2650
rect 2998 2645 3002 2649
rect 3020 2646 3027 2650
rect 3070 2645 3074 2649
rect 2849 2639 2855 2643
rect 1916 2631 1922 2635
rect 1996 2631 2000 2635
rect 2010 2631 2014 2635
rect 2028 2631 2032 2635
rect 2046 2631 2050 2635
rect 2069 2631 2073 2635
rect 2103 2631 2107 2635
rect 2118 2631 2122 2635
rect 2146 2631 2150 2635
rect 1667 2621 1671 2625
rect 1630 2615 1634 2621
rect 1646 2615 1650 2621
rect 1683 2615 1687 2621
rect 1691 2617 1695 2621
rect 1725 2621 1729 2625
rect 1928 2624 1934 2628
rect 2010 2624 2014 2628
rect 2069 2624 2073 2628
rect 2094 2624 2098 2628
rect 2125 2624 2129 2628
rect 1704 2615 1708 2621
rect 1741 2615 1745 2621
rect 2010 2616 2014 2620
rect 2053 2617 2057 2621
rect 2075 2616 2082 2620
rect 2125 2617 2129 2621
rect 1763 2612 1767 2616
rect 1996 2612 2000 2616
rect 2028 2612 2032 2616
rect 2046 2612 2050 2616
rect 2103 2612 2107 2616
rect 2118 2612 2122 2616
rect 2146 2612 2150 2616
rect 1630 2602 1634 2606
rect 1646 2602 1650 2606
rect 1691 2608 1695 2612
rect 1667 2602 1671 2608
rect 1683 2602 1687 2606
rect 1704 2602 1708 2606
rect 1725 2602 1729 2608
rect 1741 2602 1745 2606
rect 1991 2600 1995 2604
rect 1647 2589 1651 2593
rect 1691 2589 1695 2593
rect 1711 2589 1715 2593
rect 1748 2591 1752 2595
rect 2023 2598 2027 2602
rect 2043 2601 2047 2605
rect 2062 2597 2066 2601
rect 2081 2598 2085 2602
rect 2100 2598 2104 2602
rect 2113 2599 2117 2603
rect 2210 2614 2214 2618
rect 2590 2632 2594 2636
rect 2643 2632 2647 2636
rect 2693 2632 2697 2636
rect 2873 2638 2879 2642
rect 2955 2638 2959 2642
rect 3014 2638 3018 2642
rect 3039 2638 3043 2642
rect 3070 2638 3074 2642
rect 3163 2668 3167 2676
rect 3236 2690 3240 2694
rect 3190 2676 3194 2680
rect 3205 2676 3209 2680
rect 3186 2668 3190 2672
rect 3132 2662 3136 2666
rect 3145 2654 3149 2658
rect 3244 2668 3248 2676
rect 3271 2668 3275 2672
rect 3213 2662 3217 2666
rect 3226 2654 3230 2658
rect 2861 2631 2867 2635
rect 2941 2631 2945 2635
rect 2955 2631 2959 2635
rect 2973 2631 2977 2635
rect 2991 2631 2995 2635
rect 3014 2631 3018 2635
rect 3048 2631 3052 2635
rect 3063 2631 3067 2635
rect 3091 2631 3095 2635
rect 2612 2621 2616 2625
rect 2291 2614 2295 2618
rect 2575 2615 2579 2621
rect 2591 2615 2595 2621
rect 2628 2615 2632 2621
rect 2636 2617 2640 2621
rect 2670 2621 2674 2625
rect 2873 2624 2879 2628
rect 2955 2624 2959 2628
rect 3014 2624 3018 2628
rect 3039 2624 3043 2628
rect 3070 2624 3074 2628
rect 2649 2615 2653 2621
rect 2686 2615 2690 2621
rect 2955 2616 2959 2620
rect 2998 2617 3002 2621
rect 3020 2616 3027 2620
rect 3070 2617 3074 2621
rect 2708 2612 2712 2616
rect 2941 2612 2945 2616
rect 2973 2612 2977 2616
rect 2991 2612 2995 2616
rect 3048 2612 3052 2616
rect 3063 2612 3067 2616
rect 3091 2612 3095 2616
rect 2135 2598 2139 2602
rect 2143 2599 2147 2603
rect 2155 2599 2159 2603
rect 2190 2599 2194 2603
rect 2218 2598 2222 2602
rect 2270 2599 2274 2603
rect 2575 2602 2579 2606
rect 2591 2602 2595 2606
rect 2636 2608 2640 2612
rect 2612 2602 2616 2608
rect 2628 2602 2632 2606
rect 2299 2598 2303 2602
rect 2649 2602 2653 2606
rect 2670 2602 2674 2608
rect 2686 2602 2690 2606
rect 2936 2600 2940 2604
rect 1916 2582 1922 2586
rect 1996 2582 2000 2586
rect 2021 2579 2025 2583
rect 2028 2582 2032 2586
rect 2046 2582 2050 2586
rect 2068 2579 2072 2583
rect 2093 2579 2097 2583
rect 2103 2582 2107 2586
rect 2119 2582 2123 2586
rect 2139 2579 2143 2583
rect 2146 2582 2150 2586
rect 1647 2575 1651 2579
rect 1697 2575 1701 2579
rect 1748 2575 1752 2579
rect 1952 2575 1958 2579
rect 2006 2572 2010 2576
rect 2022 2572 2026 2576
rect 2053 2572 2057 2576
rect 2075 2572 2079 2576
rect 2140 2572 2144 2576
rect 2200 2578 2204 2582
rect 2592 2589 2596 2593
rect 2636 2589 2640 2593
rect 2656 2589 2660 2593
rect 2693 2591 2697 2595
rect 2968 2598 2972 2602
rect 2988 2601 2992 2605
rect 3007 2597 3011 2601
rect 3026 2598 3030 2602
rect 3045 2598 3049 2602
rect 3058 2599 3062 2603
rect 3155 2614 3159 2618
rect 3236 2614 3240 2618
rect 3080 2598 3084 2602
rect 3088 2599 3092 2603
rect 3100 2599 3104 2603
rect 3135 2599 3139 2603
rect 3163 2598 3167 2602
rect 3215 2599 3219 2603
rect 3244 2598 3248 2602
rect 2861 2582 2867 2586
rect 2941 2582 2945 2586
rect 2281 2578 2285 2582
rect 2966 2579 2970 2583
rect 2973 2582 2977 2586
rect 2991 2582 2995 2586
rect 3013 2579 3017 2583
rect 3038 2579 3042 2583
rect 3048 2582 3052 2586
rect 3064 2582 3068 2586
rect 3084 2579 3088 2583
rect 3091 2582 3095 2586
rect 2592 2575 2596 2579
rect 2642 2575 2646 2579
rect 2693 2575 2697 2579
rect 2897 2575 2903 2579
rect 2951 2572 2955 2576
rect 2967 2572 2971 2576
rect 2998 2572 3002 2576
rect 3020 2572 3024 2576
rect 3085 2572 3089 2576
rect 3145 2578 3149 2582
rect 3226 2578 3230 2582
rect 1904 2565 1910 2569
rect 1995 2565 1999 2569
rect 2029 2565 2033 2569
rect 2046 2565 2050 2569
rect 2102 2565 2106 2569
rect 2119 2565 2123 2569
rect 2147 2565 2151 2569
rect 2849 2565 2855 2569
rect 2940 2565 2944 2569
rect 2974 2565 2978 2569
rect 2991 2565 2995 2569
rect 3047 2565 3051 2569
rect 3064 2565 3068 2569
rect 3092 2565 3096 2569
rect 1940 2558 1946 2562
rect 2006 2558 2010 2562
rect 2022 2558 2026 2562
rect 2053 2558 2057 2562
rect 2075 2558 2079 2562
rect 2140 2558 2144 2562
rect 2210 2558 2214 2562
rect 1996 2548 2000 2552
rect 2021 2551 2025 2555
rect 2028 2548 2032 2552
rect 2046 2548 2050 2552
rect 2068 2551 2072 2555
rect 2093 2551 2097 2555
rect 2103 2548 2107 2552
rect 2119 2548 2123 2552
rect 2139 2551 2143 2555
rect 2146 2548 2150 2552
rect 1990 2531 1994 2535
rect 2023 2532 2027 2536
rect 2043 2529 2047 2533
rect 2062 2533 2066 2537
rect 2081 2532 2085 2536
rect 2100 2532 2104 2536
rect 2113 2531 2117 2535
rect 2135 2532 2139 2536
rect 2143 2531 2147 2535
rect 2155 2531 2159 2535
rect 2218 2536 2222 2544
rect 2315 2558 2319 2562
rect 2269 2544 2273 2548
rect 2284 2544 2288 2548
rect 2885 2558 2891 2562
rect 2951 2558 2955 2562
rect 2967 2558 2971 2562
rect 2998 2558 3002 2562
rect 3020 2558 3024 2562
rect 3085 2558 3089 2562
rect 3155 2558 3159 2562
rect 2187 2530 2191 2534
rect 2241 2535 2245 2539
rect 1996 2518 2000 2522
rect 2028 2518 2032 2522
rect 2046 2518 2050 2522
rect 2103 2518 2107 2522
rect 2118 2518 2122 2522
rect 2146 2518 2150 2522
rect 2010 2514 2014 2518
rect 2053 2513 2057 2517
rect 2075 2514 2082 2518
rect 2125 2513 2129 2517
rect 1928 2506 1934 2510
rect 2010 2506 2014 2510
rect 2069 2506 2073 2510
rect 2094 2506 2098 2510
rect 2125 2506 2129 2510
rect 2200 2522 2204 2526
rect 2323 2536 2327 2544
rect 2941 2548 2945 2552
rect 2966 2551 2970 2555
rect 2973 2548 2977 2552
rect 2991 2548 2995 2552
rect 3013 2551 3017 2555
rect 3038 2551 3042 2555
rect 3048 2548 3052 2552
rect 3064 2548 3068 2552
rect 3084 2551 3088 2555
rect 3091 2548 3095 2552
rect 2344 2536 2348 2540
rect 2292 2530 2296 2534
rect 2935 2531 2939 2535
rect 2305 2522 2309 2526
rect 2968 2532 2972 2536
rect 2988 2529 2992 2533
rect 3007 2533 3011 2537
rect 3026 2532 3030 2536
rect 3045 2532 3049 2536
rect 3058 2531 3062 2535
rect 3080 2532 3084 2536
rect 3088 2531 3092 2535
rect 3100 2531 3104 2535
rect 3163 2536 3167 2544
rect 3260 2558 3264 2562
rect 3214 2544 3218 2548
rect 3229 2544 3233 2548
rect 3132 2530 3136 2534
rect 3186 2535 3190 2539
rect 2941 2518 2945 2522
rect 2973 2518 2977 2522
rect 2991 2518 2995 2522
rect 3048 2518 3052 2522
rect 3063 2518 3067 2522
rect 3091 2518 3095 2522
rect 2955 2514 2959 2518
rect 2998 2513 3002 2517
rect 3020 2514 3027 2518
rect 3070 2513 3074 2517
rect 2873 2506 2879 2510
rect 2955 2506 2959 2510
rect 3014 2506 3018 2510
rect 3039 2506 3043 2510
rect 3070 2506 3074 2510
rect 3145 2522 3149 2526
rect 3268 2536 3272 2544
rect 3289 2536 3293 2540
rect 3237 2530 3241 2534
rect 3250 2522 3254 2526
rect 1916 2499 1922 2503
rect 1996 2499 2000 2503
rect 2010 2499 2014 2503
rect 2028 2499 2032 2503
rect 2046 2499 2050 2503
rect 2069 2499 2073 2503
rect 2103 2499 2107 2503
rect 2118 2499 2122 2503
rect 2146 2499 2150 2503
rect 2861 2499 2867 2503
rect 2941 2499 2945 2503
rect 2955 2499 2959 2503
rect 2973 2499 2977 2503
rect 2991 2499 2995 2503
rect 3014 2499 3018 2503
rect 3048 2499 3052 2503
rect 3063 2499 3067 2503
rect 3091 2499 3095 2503
rect 1928 2492 1934 2496
rect 2010 2492 2014 2496
rect 2069 2492 2073 2496
rect 2094 2492 2098 2496
rect 2125 2492 2129 2496
rect 2010 2484 2014 2488
rect 2053 2485 2057 2489
rect 2075 2484 2082 2488
rect 2125 2485 2129 2489
rect 1996 2480 2000 2484
rect 2028 2480 2032 2484
rect 2046 2480 2050 2484
rect 2103 2480 2107 2484
rect 2118 2480 2122 2484
rect 2146 2480 2150 2484
rect 2210 2483 2214 2487
rect 2873 2492 2879 2496
rect 2955 2492 2959 2496
rect 3014 2492 3018 2496
rect 3039 2492 3043 2496
rect 3070 2492 3074 2496
rect 2315 2483 2319 2487
rect 2955 2484 2959 2488
rect 2998 2485 3002 2489
rect 3020 2484 3027 2488
rect 3070 2485 3074 2489
rect 2941 2480 2945 2484
rect 2973 2480 2977 2484
rect 2991 2480 2995 2484
rect 3048 2480 3052 2484
rect 3063 2480 3067 2484
rect 3091 2480 3095 2484
rect 3155 2483 3159 2487
rect 3260 2483 3264 2487
rect 1991 2468 1995 2472
rect 2023 2466 2027 2470
rect 2043 2469 2047 2473
rect 2062 2465 2066 2469
rect 2081 2466 2085 2470
rect 2100 2466 2104 2470
rect 2113 2467 2117 2471
rect 2135 2466 2139 2470
rect 2143 2467 2147 2471
rect 2155 2467 2159 2471
rect 2189 2468 2193 2472
rect 2218 2467 2222 2471
rect 2295 2468 2299 2472
rect 2323 2467 2327 2471
rect 2936 2468 2940 2472
rect 1996 2450 2000 2454
rect 2021 2447 2025 2451
rect 2028 2450 2032 2454
rect 2046 2450 2050 2454
rect 2068 2447 2072 2451
rect 2093 2447 2097 2451
rect 2103 2450 2107 2454
rect 2119 2450 2123 2454
rect 2139 2447 2143 2451
rect 2146 2450 2150 2454
rect 1940 2440 1946 2444
rect 2022 2440 2026 2444
rect 2053 2440 2057 2444
rect 2075 2440 2079 2444
rect 2140 2440 2144 2444
rect 2200 2447 2204 2451
rect 2968 2466 2972 2470
rect 2988 2469 2992 2473
rect 3007 2465 3011 2469
rect 3026 2466 3030 2470
rect 3045 2466 3049 2470
rect 3058 2467 3062 2471
rect 3080 2466 3084 2470
rect 3088 2467 3092 2471
rect 3100 2467 3104 2471
rect 3134 2468 3138 2472
rect 3163 2467 3167 2471
rect 3240 2468 3244 2472
rect 3268 2467 3272 2471
rect 2305 2447 2309 2451
rect 2941 2450 2945 2454
rect 2966 2447 2970 2451
rect 2973 2450 2977 2454
rect 2991 2450 2995 2454
rect 3013 2447 3017 2451
rect 3038 2447 3042 2451
rect 3048 2450 3052 2454
rect 3064 2450 3068 2454
rect 3084 2447 3088 2451
rect 3091 2450 3095 2454
rect 2885 2440 2891 2444
rect 2967 2440 2971 2444
rect 2998 2440 3002 2444
rect 3020 2440 3024 2444
rect 3085 2440 3089 2444
rect 3145 2447 3149 2451
rect 3250 2447 3254 2451
rect 1904 2433 1910 2437
rect 1995 2433 1999 2437
rect 2029 2433 2033 2437
rect 2046 2433 2050 2437
rect 2102 2433 2106 2437
rect 2119 2433 2123 2437
rect 2147 2433 2151 2437
rect 2849 2433 2855 2437
rect 2940 2433 2944 2437
rect 2974 2433 2978 2437
rect 2991 2433 2995 2437
rect 3047 2433 3051 2437
rect 3064 2433 3068 2437
rect 3092 2433 3096 2437
rect 1940 2426 1946 2430
rect 2022 2426 2026 2430
rect 2053 2426 2057 2430
rect 2075 2426 2079 2430
rect 2140 2426 2144 2430
rect 2210 2426 2214 2430
rect 1996 2416 2000 2420
rect 2021 2419 2025 2423
rect 2028 2416 2032 2420
rect 2046 2416 2050 2420
rect 2068 2419 2072 2423
rect 2093 2419 2097 2423
rect 2103 2416 2107 2420
rect 2119 2416 2123 2420
rect 2139 2419 2143 2423
rect 2146 2416 2150 2420
rect 1990 2399 1994 2403
rect 2023 2400 2027 2404
rect 2043 2397 2047 2401
rect 2062 2401 2066 2405
rect 2081 2400 2085 2404
rect 2100 2400 2104 2404
rect 2113 2399 2117 2403
rect 2135 2400 2139 2404
rect 2143 2399 2147 2403
rect 2155 2399 2159 2403
rect 2218 2404 2222 2412
rect 2291 2426 2295 2430
rect 2245 2412 2249 2416
rect 2260 2412 2264 2416
rect 2241 2404 2245 2408
rect 2187 2398 2191 2402
rect 1996 2386 2000 2390
rect 2028 2386 2032 2390
rect 2046 2386 2050 2390
rect 2103 2386 2107 2390
rect 2118 2386 2122 2390
rect 2146 2386 2150 2390
rect 2010 2382 2014 2386
rect 2053 2381 2057 2385
rect 2075 2382 2082 2386
rect 2125 2381 2129 2385
rect 1928 2374 1934 2378
rect 2010 2374 2014 2378
rect 2069 2374 2073 2378
rect 2094 2374 2098 2378
rect 2125 2374 2129 2378
rect 2200 2390 2204 2394
rect 2299 2404 2303 2412
rect 2381 2426 2385 2430
rect 2335 2412 2339 2416
rect 2350 2412 2354 2416
rect 2885 2426 2891 2430
rect 2967 2426 2971 2430
rect 2998 2426 3002 2430
rect 3020 2426 3024 2430
rect 3085 2426 3089 2430
rect 3155 2426 3159 2430
rect 2323 2404 2327 2408
rect 2268 2398 2272 2402
rect 2357 2406 2361 2410
rect 2389 2404 2393 2412
rect 2941 2416 2945 2420
rect 2966 2419 2970 2423
rect 2973 2416 2977 2420
rect 2991 2416 2995 2420
rect 3013 2419 3017 2423
rect 3038 2419 3042 2423
rect 3048 2416 3052 2420
rect 3064 2416 3068 2420
rect 3084 2419 3088 2423
rect 3091 2416 3095 2420
rect 2281 2390 2285 2394
rect 2424 2403 2428 2407
rect 2935 2399 2939 2403
rect 2371 2390 2375 2394
rect 2968 2400 2972 2404
rect 2988 2397 2992 2401
rect 3007 2401 3011 2405
rect 3026 2400 3030 2404
rect 3045 2400 3049 2404
rect 3058 2399 3062 2403
rect 3080 2400 3084 2404
rect 3088 2399 3092 2403
rect 3100 2399 3104 2403
rect 3163 2404 3167 2412
rect 3236 2426 3240 2430
rect 3190 2412 3194 2416
rect 3205 2412 3209 2416
rect 3186 2404 3190 2408
rect 3132 2398 3136 2402
rect 2941 2386 2945 2390
rect 2973 2386 2977 2390
rect 2991 2386 2995 2390
rect 3048 2386 3052 2390
rect 3063 2386 3067 2390
rect 3091 2386 3095 2390
rect 2955 2382 2959 2386
rect 2998 2381 3002 2385
rect 3020 2382 3027 2386
rect 3070 2381 3074 2385
rect 2873 2374 2879 2378
rect 2955 2374 2959 2378
rect 3014 2374 3018 2378
rect 3039 2374 3043 2378
rect 3070 2374 3074 2378
rect 3145 2390 3149 2394
rect 3244 2404 3248 2412
rect 3326 2426 3330 2430
rect 3280 2412 3284 2416
rect 3295 2412 3299 2416
rect 3268 2404 3272 2408
rect 3213 2398 3217 2402
rect 3302 2406 3306 2410
rect 3334 2404 3338 2412
rect 3226 2390 3230 2394
rect 3369 2403 3373 2407
rect 4228 2403 4240 2407
rect 3316 2390 3320 2394
rect 1916 2367 1922 2371
rect 1996 2367 2000 2371
rect 2010 2367 2014 2371
rect 2028 2367 2032 2371
rect 2046 2367 2050 2371
rect 2069 2367 2073 2371
rect 2103 2367 2107 2371
rect 2118 2367 2122 2371
rect 2146 2367 2150 2371
rect 2861 2367 2867 2371
rect 2941 2367 2945 2371
rect 2955 2367 2959 2371
rect 2973 2367 2977 2371
rect 2991 2367 2995 2371
rect 3014 2367 3018 2371
rect 3048 2367 3052 2371
rect 3063 2367 3067 2371
rect 3091 2367 3095 2371
rect 1928 2360 1934 2364
rect 2010 2360 2014 2364
rect 2069 2360 2073 2364
rect 2094 2360 2098 2364
rect 2125 2360 2129 2364
rect 2010 2352 2014 2356
rect 2053 2353 2057 2357
rect 2075 2352 2082 2356
rect 2125 2353 2129 2357
rect 1996 2348 2000 2352
rect 2028 2348 2032 2352
rect 2046 2348 2050 2352
rect 2103 2348 2107 2352
rect 2118 2348 2122 2352
rect 2146 2348 2150 2352
rect 1991 2336 1995 2340
rect 2023 2334 2027 2338
rect 2043 2337 2047 2341
rect 2062 2333 2066 2337
rect 2081 2334 2085 2338
rect 2100 2334 2104 2338
rect 2113 2335 2117 2339
rect 2210 2348 2214 2352
rect 2291 2348 2295 2352
rect 2873 2360 2879 2364
rect 2955 2360 2959 2364
rect 3014 2360 3018 2364
rect 3039 2360 3043 2364
rect 3070 2360 3074 2364
rect 2955 2352 2959 2356
rect 2998 2353 3002 2357
rect 3020 2352 3027 2356
rect 3070 2353 3074 2357
rect 2381 2348 2385 2352
rect 2941 2348 2945 2352
rect 2973 2348 2977 2352
rect 2991 2348 2995 2352
rect 3048 2348 3052 2352
rect 3063 2348 3067 2352
rect 3091 2348 3095 2352
rect 2135 2334 2139 2338
rect 2143 2335 2147 2339
rect 2155 2335 2159 2339
rect 2190 2333 2194 2337
rect 2218 2332 2222 2336
rect 2270 2333 2274 2337
rect 2299 2332 2303 2336
rect 2354 2333 2358 2337
rect 2936 2336 2940 2340
rect 2389 2332 2393 2336
rect 1996 2318 2000 2322
rect 2021 2315 2025 2319
rect 2028 2318 2032 2322
rect 2046 2318 2050 2322
rect 2068 2315 2072 2319
rect 2093 2315 2097 2319
rect 2103 2318 2107 2322
rect 2119 2318 2123 2322
rect 2139 2315 2143 2319
rect 2146 2318 2150 2322
rect 2968 2334 2972 2338
rect 2988 2337 2992 2341
rect 3007 2333 3011 2337
rect 3026 2334 3030 2338
rect 3045 2334 3049 2338
rect 3058 2335 3062 2339
rect 3155 2348 3159 2352
rect 3236 2348 3240 2352
rect 3326 2348 3330 2352
rect 4228 2342 4240 2355
rect 3080 2334 3084 2338
rect 3088 2335 3092 2339
rect 3100 2335 3104 2339
rect 3135 2333 3139 2337
rect 3163 2332 3167 2336
rect 3215 2333 3219 2337
rect 3244 2332 3248 2336
rect 3299 2333 3303 2337
rect 3334 2332 3338 2336
rect 1940 2308 1946 2312
rect 2022 2308 2026 2312
rect 2053 2308 2057 2312
rect 2075 2308 2079 2312
rect 2140 2308 2144 2312
rect 2200 2312 2204 2316
rect 2281 2312 2285 2316
rect 2941 2318 2945 2322
rect 2371 2312 2375 2316
rect 2966 2315 2970 2319
rect 2973 2318 2977 2322
rect 2991 2318 2995 2322
rect 3013 2315 3017 2319
rect 3038 2315 3042 2319
rect 3048 2318 3052 2322
rect 3064 2318 3068 2322
rect 3084 2315 3088 2319
rect 3091 2318 3095 2322
rect 2885 2308 2891 2312
rect 2967 2308 2971 2312
rect 2998 2308 3002 2312
rect 3020 2308 3024 2312
rect 3085 2308 3089 2312
rect 3145 2312 3149 2316
rect 3226 2312 3230 2316
rect 3316 2312 3320 2316
rect 1904 2301 1910 2305
rect 1995 2301 1999 2305
rect 2029 2301 2033 2305
rect 2046 2301 2050 2305
rect 2102 2301 2106 2305
rect 2119 2301 2123 2305
rect 2147 2301 2151 2305
rect 2849 2301 2855 2305
rect 2940 2301 2944 2305
rect 2974 2301 2978 2305
rect 2991 2301 2995 2305
rect 3047 2301 3051 2305
rect 3064 2301 3068 2305
rect 3092 2301 3096 2305
rect 1940 2294 1946 2298
rect 2022 2294 2026 2298
rect 2053 2294 2057 2298
rect 2075 2294 2079 2298
rect 2140 2294 2144 2298
rect 2210 2294 2214 2298
rect 1996 2284 2000 2288
rect 2021 2287 2025 2291
rect 2028 2284 2032 2288
rect 2046 2284 2050 2288
rect 2068 2287 2072 2291
rect 2093 2287 2097 2291
rect 2103 2284 2107 2288
rect 2119 2284 2123 2288
rect 2139 2287 2143 2291
rect 2146 2284 2150 2288
rect 1990 2267 1994 2271
rect 2023 2268 2027 2272
rect 2043 2265 2047 2269
rect 2062 2269 2066 2273
rect 2885 2294 2891 2298
rect 2967 2294 2971 2298
rect 2998 2294 3002 2298
rect 3020 2294 3024 2298
rect 3085 2294 3089 2298
rect 3155 2294 3159 2298
rect 2081 2268 2085 2272
rect 2100 2268 2104 2272
rect 2113 2267 2117 2271
rect 2135 2268 2139 2272
rect 2143 2267 2147 2271
rect 2155 2267 2159 2271
rect 2218 2272 2222 2280
rect 2941 2284 2945 2288
rect 2966 2287 2970 2291
rect 2973 2284 2977 2288
rect 2991 2284 2995 2288
rect 3013 2287 3017 2291
rect 3038 2287 3042 2291
rect 3048 2284 3052 2288
rect 3064 2284 3068 2288
rect 3084 2287 3088 2291
rect 3091 2284 3095 2288
rect 2187 2266 2191 2270
rect 2241 2271 2245 2275
rect 2935 2267 2939 2271
rect 1996 2254 2000 2258
rect 2028 2254 2032 2258
rect 2046 2254 2050 2258
rect 2103 2254 2107 2258
rect 2118 2254 2122 2258
rect 2146 2254 2150 2258
rect 2010 2250 2014 2254
rect 1513 2246 1517 2250
rect 1549 2246 1553 2250
rect 1616 2246 1620 2250
rect 1645 2246 1649 2250
rect 1681 2246 1685 2250
rect 1748 2246 1752 2250
rect 1777 2246 1781 2250
rect 1813 2246 1817 2250
rect 1880 2246 1884 2250
rect 1964 2246 1970 2250
rect 2053 2249 2057 2253
rect 2075 2250 2082 2254
rect 2125 2249 2129 2253
rect 1904 2239 1910 2243
rect 2010 2242 2014 2246
rect 2019 2242 2023 2246
rect 2069 2242 2073 2246
rect 2094 2242 2098 2246
rect 2125 2242 2129 2246
rect 2200 2258 2204 2262
rect 2968 2268 2972 2272
rect 2988 2265 2992 2269
rect 3007 2269 3011 2273
rect 3026 2268 3030 2272
rect 3045 2268 3049 2272
rect 3058 2267 3062 2271
rect 3080 2268 3084 2272
rect 3088 2267 3092 2271
rect 3100 2267 3104 2271
rect 3163 2272 3167 2280
rect 3132 2266 3136 2270
rect 3186 2271 3190 2275
rect 2941 2254 2945 2258
rect 2973 2254 2977 2258
rect 2991 2254 2995 2258
rect 3048 2254 3052 2258
rect 3063 2254 3067 2258
rect 3091 2254 3095 2258
rect 2955 2250 2959 2254
rect 2458 2246 2462 2250
rect 2494 2246 2498 2250
rect 2561 2246 2565 2250
rect 2590 2246 2594 2250
rect 2626 2246 2630 2250
rect 2693 2246 2697 2250
rect 2722 2246 2726 2250
rect 2758 2246 2762 2250
rect 2825 2246 2829 2250
rect 2909 2246 2915 2250
rect 2998 2249 3002 2253
rect 3020 2250 3027 2254
rect 3070 2249 3074 2253
rect 2849 2239 2855 2243
rect 2955 2242 2959 2246
rect 2964 2242 2968 2246
rect 3014 2242 3018 2246
rect 3039 2242 3043 2246
rect 3070 2242 3074 2246
rect 3145 2258 3149 2262
rect 1513 2232 1517 2236
rect 1563 2232 1567 2236
rect 1616 2232 1620 2236
rect 1645 2232 1649 2236
rect 1695 2232 1699 2236
rect 1748 2232 1752 2236
rect 1777 2232 1781 2236
rect 1827 2232 1831 2236
rect 1880 2232 1884 2236
rect 1916 2235 1922 2239
rect 1996 2235 2000 2239
rect 2010 2235 2014 2239
rect 2028 2235 2032 2239
rect 2046 2235 2050 2239
rect 2069 2235 2073 2239
rect 2103 2235 2107 2239
rect 2118 2235 2122 2239
rect 2146 2235 2150 2239
rect 2271 2235 2275 2239
rect 2289 2235 2293 2239
rect 2307 2235 2311 2239
rect 2330 2235 2334 2239
rect 2364 2235 2368 2239
rect 2379 2235 2383 2239
rect 2407 2235 2411 2239
rect 1536 2221 1540 2225
rect 1507 2212 1511 2216
rect 1520 2215 1524 2221
rect 1557 2215 1561 2221
rect 1570 2217 1574 2221
rect 1594 2221 1598 2225
rect 1668 2221 1672 2225
rect 1578 2215 1582 2221
rect 1615 2215 1619 2221
rect 1631 2215 1635 2221
rect 1652 2215 1656 2221
rect 1689 2215 1693 2221
rect 1702 2217 1706 2221
rect 1726 2221 1730 2225
rect 1800 2221 1804 2225
rect 1710 2215 1714 2221
rect 1747 2215 1751 2221
rect 1763 2215 1767 2221
rect 1784 2215 1788 2221
rect 1821 2215 1825 2221
rect 1834 2217 1838 2221
rect 1858 2221 1862 2225
rect 1928 2228 1934 2232
rect 2010 2228 2014 2232
rect 2019 2228 2023 2232
rect 2069 2228 2073 2232
rect 2094 2228 2098 2232
rect 2125 2228 2129 2232
rect 1842 2215 1846 2221
rect 1879 2215 1883 2221
rect 1895 2217 1899 2221
rect 2010 2220 2014 2224
rect 2053 2221 2057 2225
rect 2075 2220 2082 2224
rect 2125 2221 2129 2225
rect 1996 2216 2000 2220
rect 2028 2216 2032 2220
rect 2046 2216 2050 2220
rect 2103 2216 2107 2220
rect 2118 2216 2122 2220
rect 2146 2216 2150 2220
rect 1520 2202 1524 2206
rect 1536 2202 1540 2208
rect 1570 2208 1574 2212
rect 1557 2202 1561 2206
rect 1578 2202 1582 2206
rect 1594 2202 1598 2208
rect 1615 2202 1619 2206
rect 1631 2202 1635 2206
rect 1652 2202 1656 2206
rect 1668 2202 1672 2208
rect 1702 2208 1706 2212
rect 1689 2202 1693 2206
rect 1710 2202 1714 2206
rect 1726 2202 1730 2208
rect 1747 2202 1751 2206
rect 1763 2202 1767 2206
rect 1784 2202 1788 2206
rect 1800 2202 1804 2208
rect 1834 2208 1838 2212
rect 1821 2202 1825 2206
rect 1842 2202 1846 2206
rect 1858 2202 1862 2208
rect 1879 2202 1883 2206
rect 1895 2202 1899 2206
rect 1991 2204 1995 2208
rect 1513 2191 1517 2195
rect 1550 2189 1554 2193
rect 1570 2189 1574 2193
rect 1614 2189 1618 2193
rect 1645 2191 1649 2195
rect 1682 2189 1686 2193
rect 1702 2189 1706 2193
rect 1746 2189 1750 2193
rect 1777 2191 1781 2195
rect 1814 2189 1818 2193
rect 1834 2189 1838 2193
rect 1878 2189 1882 2193
rect 2023 2202 2027 2206
rect 2043 2205 2047 2209
rect 2062 2201 2066 2205
rect 2081 2202 2085 2206
rect 2100 2202 2104 2206
rect 2113 2203 2117 2207
rect 2249 2228 2253 2232
rect 2271 2228 2275 2232
rect 2330 2228 2334 2232
rect 2355 2228 2359 2232
rect 2386 2228 2390 2232
rect 2458 2232 2462 2236
rect 2508 2232 2512 2236
rect 2561 2232 2565 2236
rect 2590 2232 2594 2236
rect 2640 2232 2644 2236
rect 2693 2232 2697 2236
rect 2722 2232 2726 2236
rect 2772 2232 2776 2236
rect 2825 2232 2829 2236
rect 2861 2235 2867 2239
rect 2941 2235 2945 2239
rect 2955 2235 2959 2239
rect 2973 2235 2977 2239
rect 2991 2235 2995 2239
rect 3014 2235 3018 2239
rect 3048 2235 3052 2239
rect 3063 2235 3067 2239
rect 3091 2235 3095 2239
rect 3216 2235 3220 2239
rect 3234 2235 3238 2239
rect 3252 2235 3256 2239
rect 3275 2235 3279 2239
rect 3309 2235 3313 2239
rect 3324 2235 3328 2239
rect 3352 2235 3356 2239
rect 2271 2220 2275 2224
rect 2314 2221 2318 2225
rect 2336 2220 2343 2224
rect 2386 2221 2390 2225
rect 2481 2221 2485 2225
rect 2289 2216 2293 2220
rect 2307 2216 2311 2220
rect 2364 2216 2368 2220
rect 2379 2216 2383 2220
rect 2407 2216 2411 2220
rect 2210 2212 2214 2216
rect 2135 2202 2139 2206
rect 2143 2203 2147 2207
rect 2155 2203 2159 2207
rect 2189 2197 2193 2201
rect 2229 2203 2233 2207
rect 2218 2196 2222 2200
rect 1996 2186 2000 2190
rect 1916 2182 1922 2186
rect 2021 2183 2025 2187
rect 2028 2186 2032 2190
rect 2046 2186 2050 2190
rect 2068 2183 2072 2187
rect 2093 2183 2097 2187
rect 2103 2186 2107 2190
rect 2119 2186 2123 2190
rect 2139 2183 2143 2187
rect 2146 2186 2150 2190
rect 2284 2202 2288 2206
rect 2304 2205 2308 2209
rect 2323 2201 2327 2205
rect 2452 2212 2456 2216
rect 2465 2215 2469 2221
rect 2502 2215 2506 2221
rect 2515 2217 2519 2221
rect 2539 2221 2543 2225
rect 2613 2221 2617 2225
rect 2523 2215 2527 2221
rect 2560 2215 2564 2221
rect 2576 2215 2580 2221
rect 2597 2215 2601 2221
rect 2634 2215 2638 2221
rect 2647 2217 2651 2221
rect 2671 2221 2675 2225
rect 2745 2221 2749 2225
rect 2655 2215 2659 2221
rect 2692 2215 2696 2221
rect 2708 2215 2712 2221
rect 2729 2215 2733 2221
rect 2766 2215 2770 2221
rect 2779 2217 2783 2221
rect 2803 2221 2807 2225
rect 2873 2228 2879 2232
rect 2955 2228 2959 2232
rect 2964 2228 2968 2232
rect 3014 2228 3018 2232
rect 3039 2228 3043 2232
rect 3070 2228 3074 2232
rect 2787 2215 2791 2221
rect 2824 2215 2828 2221
rect 2840 2217 2844 2221
rect 2955 2220 2959 2224
rect 2998 2221 3002 2225
rect 3020 2220 3027 2224
rect 3070 2221 3074 2225
rect 2941 2216 2945 2220
rect 2973 2216 2977 2220
rect 2991 2216 2995 2220
rect 3048 2216 3052 2220
rect 3063 2216 3067 2220
rect 3091 2216 3095 2220
rect 2342 2202 2346 2206
rect 2361 2202 2365 2206
rect 2374 2203 2378 2207
rect 2396 2202 2400 2206
rect 2404 2203 2408 2207
rect 2416 2203 2420 2207
rect 2465 2202 2469 2206
rect 2481 2202 2485 2208
rect 2515 2208 2519 2212
rect 2502 2202 2506 2206
rect 2523 2202 2527 2206
rect 2539 2202 2543 2208
rect 2560 2202 2564 2206
rect 2576 2202 2580 2206
rect 2597 2202 2601 2206
rect 2613 2202 2617 2208
rect 2647 2208 2651 2212
rect 2634 2202 2638 2206
rect 2655 2202 2659 2206
rect 2671 2202 2675 2208
rect 2692 2202 2696 2206
rect 2708 2202 2712 2206
rect 2729 2202 2733 2206
rect 2745 2202 2749 2208
rect 2779 2208 2783 2212
rect 2766 2202 2770 2206
rect 2787 2202 2791 2206
rect 2803 2202 2807 2208
rect 2824 2202 2828 2206
rect 2840 2202 2844 2206
rect 2936 2204 2940 2208
rect 2230 2186 2234 2190
rect 2256 2186 2260 2190
rect 1513 2175 1517 2179
rect 1564 2175 1568 2179
rect 1614 2175 1618 2179
rect 1645 2175 1649 2179
rect 1696 2175 1700 2179
rect 1746 2175 1750 2179
rect 1777 2175 1781 2179
rect 1828 2175 1832 2179
rect 1878 2175 1882 2179
rect 1952 2176 1958 2180
rect 2004 2176 2008 2180
rect 2022 2176 2026 2180
rect 2053 2176 2057 2180
rect 2075 2176 2079 2180
rect 2140 2176 2144 2180
rect 2282 2183 2286 2187
rect 2289 2186 2293 2190
rect 2307 2186 2311 2190
rect 2329 2183 2333 2187
rect 2354 2183 2358 2187
rect 2364 2186 2368 2190
rect 2380 2186 2384 2190
rect 2400 2183 2404 2187
rect 2407 2186 2411 2190
rect 2458 2191 2462 2195
rect 2495 2189 2499 2193
rect 2515 2189 2519 2193
rect 2559 2189 2563 2193
rect 2590 2191 2594 2195
rect 2627 2189 2631 2193
rect 2647 2189 2651 2193
rect 2691 2189 2695 2193
rect 2722 2191 2726 2195
rect 2759 2189 2763 2193
rect 2779 2189 2783 2193
rect 2823 2189 2827 2193
rect 2968 2202 2972 2206
rect 2988 2205 2992 2209
rect 3007 2201 3011 2205
rect 3026 2202 3030 2206
rect 3045 2202 3049 2206
rect 3058 2203 3062 2207
rect 3194 2228 3198 2232
rect 3216 2228 3220 2232
rect 3275 2228 3279 2232
rect 3300 2228 3304 2232
rect 3331 2228 3335 2232
rect 3216 2220 3220 2224
rect 3259 2221 3263 2225
rect 3281 2220 3288 2224
rect 3331 2221 3335 2225
rect 3234 2216 3238 2220
rect 3252 2216 3256 2220
rect 3309 2216 3313 2220
rect 3324 2216 3328 2220
rect 3352 2216 3356 2220
rect 3155 2212 3159 2216
rect 3080 2202 3084 2206
rect 3088 2203 3092 2207
rect 3100 2203 3104 2207
rect 3134 2197 3138 2201
rect 3174 2203 3178 2207
rect 3163 2196 3167 2200
rect 2941 2186 2945 2190
rect 2861 2182 2867 2186
rect 2966 2183 2970 2187
rect 2973 2186 2977 2190
rect 2991 2186 2995 2190
rect 3013 2183 3017 2187
rect 3038 2183 3042 2187
rect 3048 2186 3052 2190
rect 3064 2186 3068 2190
rect 3084 2183 3088 2187
rect 3091 2186 3095 2190
rect 3229 2202 3233 2206
rect 3249 2205 3253 2209
rect 3268 2201 3272 2205
rect 3287 2202 3291 2206
rect 3306 2202 3310 2206
rect 3319 2203 3323 2207
rect 3341 2202 3345 2206
rect 3349 2203 3353 2207
rect 3361 2203 3365 2207
rect 3175 2186 3179 2190
rect 3201 2186 3205 2190
rect 2200 2176 2204 2180
rect 2239 2176 2243 2180
rect 2283 2176 2287 2180
rect 2314 2176 2318 2180
rect 2336 2176 2340 2180
rect 2401 2176 2405 2180
rect 2458 2175 2462 2179
rect 2509 2175 2513 2179
rect 2559 2175 2563 2179
rect 2590 2175 2594 2179
rect 2641 2175 2645 2179
rect 2691 2175 2695 2179
rect 2722 2175 2726 2179
rect 2773 2175 2777 2179
rect 2823 2175 2827 2179
rect 2897 2176 2903 2180
rect 2949 2176 2953 2180
rect 2967 2176 2971 2180
rect 2998 2176 3002 2180
rect 3020 2176 3024 2180
rect 3085 2176 3089 2180
rect 3227 2183 3231 2187
rect 3234 2186 3238 2190
rect 3252 2186 3256 2190
rect 3274 2183 3278 2187
rect 3299 2183 3303 2187
rect 3309 2186 3313 2190
rect 3325 2186 3329 2190
rect 3345 2183 3349 2187
rect 3352 2186 3356 2190
rect 3145 2176 3149 2180
rect 3184 2176 3188 2180
rect 3228 2176 3232 2180
rect 3259 2176 3263 2180
rect 3281 2176 3285 2180
rect 3346 2176 3350 2180
rect 1507 2168 1511 2172
rect 1895 2168 1899 2172
rect 1904 2169 1910 2173
rect 1995 2169 1999 2173
rect 2029 2169 2033 2173
rect 2046 2169 2050 2173
rect 2102 2169 2106 2173
rect 2119 2169 2123 2173
rect 2147 2169 2151 2173
rect 2230 2169 2234 2173
rect 2256 2169 2260 2173
rect 2290 2169 2294 2173
rect 2307 2169 2311 2173
rect 2363 2169 2367 2173
rect 2380 2169 2384 2173
rect 2408 2169 2412 2173
rect 2452 2168 2456 2172
rect 2840 2168 2844 2172
rect 2849 2169 2855 2173
rect 2940 2169 2944 2173
rect 2974 2169 2978 2173
rect 2991 2169 2995 2173
rect 3047 2169 3051 2173
rect 3064 2169 3068 2173
rect 3092 2169 3096 2173
rect 3175 2169 3179 2173
rect 3201 2169 3205 2173
rect 3235 2169 3239 2173
rect 3252 2169 3256 2173
rect 3308 2169 3312 2173
rect 3325 2169 3329 2173
rect 3353 2169 3357 2173
rect 1630 2161 1635 2165
rect 1763 2161 1767 2165
rect 1940 2162 1946 2166
rect 2004 2162 2008 2166
rect 2238 2162 2242 2166
rect 2424 2163 2428 2167
rect 2436 2163 2440 2167
rect 2575 2161 2580 2165
rect 2708 2161 2712 2165
rect 2885 2162 2891 2166
rect 2949 2162 2953 2166
rect 3183 2162 3187 2166
rect 3369 2163 3373 2167
rect 3381 2163 3385 2167
rect 1638 2154 1642 2158
rect 1928 2154 1934 2158
rect 2248 2155 2252 2159
rect 2413 2155 2417 2159
rect 1622 2150 1626 2154
rect 1654 2150 1658 2154
rect 1976 2148 1982 2152
rect 2583 2154 2587 2158
rect 2873 2154 2879 2158
rect 3193 2155 3197 2159
rect 3358 2155 3362 2159
rect 2567 2150 2571 2154
rect 2599 2150 2603 2154
rect 2921 2148 2927 2152
rect 1622 2141 1626 2145
rect 1654 2141 1658 2145
rect 2567 2141 2571 2145
rect 2599 2141 2603 2145
rect 1638 2134 1642 2138
rect 1895 2134 1899 2138
rect 1964 2134 1970 2138
rect 2296 2134 2300 2138
rect 2332 2134 2336 2138
rect 2399 2134 2403 2138
rect 2583 2134 2587 2138
rect 2840 2134 2844 2138
rect 2909 2134 2915 2138
rect 3241 2134 3245 2138
rect 3277 2134 3281 2138
rect 3344 2134 3348 2138
rect 1895 2126 1899 2130
rect 1904 2127 1910 2131
rect 2282 2127 2286 2131
rect 1622 2122 1626 2126
rect 1654 2122 1658 2126
rect 1638 2118 1642 2122
rect 2296 2120 2300 2124
rect 2346 2120 2350 2124
rect 2399 2120 2403 2124
rect 2840 2126 2844 2130
rect 2849 2127 2855 2131
rect 3227 2127 3231 2131
rect 2567 2122 2571 2126
rect 2599 2122 2603 2126
rect 2583 2118 2587 2122
rect 3241 2120 3245 2124
rect 3291 2120 3295 2124
rect 3344 2120 3348 2124
rect 1630 2111 1635 2115
rect 1764 2111 1768 2115
rect 2319 2109 2323 2113
rect 1513 2104 1517 2108
rect 1549 2104 1553 2108
rect 1616 2104 1620 2108
rect 1645 2104 1649 2108
rect 1681 2104 1685 2108
rect 1748 2104 1752 2108
rect 1777 2104 1781 2108
rect 1813 2104 1817 2108
rect 1880 2104 1884 2108
rect 1964 2104 1970 2108
rect 1904 2097 1910 2101
rect 2290 2100 2294 2104
rect 2303 2103 2307 2109
rect 2340 2103 2344 2109
rect 2353 2105 2357 2109
rect 2377 2109 2381 2113
rect 2575 2111 2580 2115
rect 2709 2111 2713 2115
rect 3264 2109 3268 2113
rect 2361 2103 2365 2109
rect 2398 2103 2402 2109
rect 2414 2103 2418 2109
rect 2458 2104 2462 2108
rect 2494 2104 2498 2108
rect 2561 2104 2565 2108
rect 2590 2104 2594 2108
rect 2626 2104 2630 2108
rect 2693 2104 2697 2108
rect 2722 2104 2726 2108
rect 2758 2104 2762 2108
rect 2825 2104 2829 2108
rect 2909 2104 2915 2108
rect 1513 2090 1517 2094
rect 1563 2090 1567 2094
rect 1616 2090 1620 2094
rect 1645 2090 1649 2094
rect 1695 2090 1699 2094
rect 1748 2090 1752 2094
rect 1777 2090 1781 2094
rect 1827 2090 1831 2094
rect 1880 2090 1884 2094
rect 2303 2090 2307 2094
rect 2319 2090 2323 2096
rect 2353 2096 2357 2100
rect 2340 2090 2344 2094
rect 1536 2079 1540 2083
rect 1507 2070 1511 2074
rect 1520 2073 1524 2079
rect 1557 2073 1561 2079
rect 1570 2075 1574 2079
rect 1594 2079 1598 2083
rect 1668 2079 1672 2083
rect 1578 2073 1582 2079
rect 1615 2073 1619 2079
rect 1631 2073 1635 2079
rect 1652 2073 1656 2079
rect 1689 2073 1693 2079
rect 1702 2075 1706 2079
rect 1726 2079 1730 2083
rect 1800 2079 1804 2083
rect 1710 2073 1714 2079
rect 1747 2073 1751 2079
rect 1763 2073 1767 2079
rect 1784 2073 1788 2079
rect 1821 2073 1825 2079
rect 1834 2075 1838 2079
rect 1858 2079 1862 2083
rect 1842 2073 1846 2079
rect 1879 2073 1883 2079
rect 1895 2075 1899 2079
rect 2361 2090 2365 2094
rect 2377 2090 2381 2096
rect 2849 2097 2855 2101
rect 3235 2100 3239 2104
rect 3248 2103 3252 2109
rect 3285 2103 3289 2109
rect 3298 2105 3302 2109
rect 3322 2109 3326 2113
rect 3306 2103 3310 2109
rect 3343 2103 3347 2109
rect 3359 2103 3363 2109
rect 2398 2090 2402 2094
rect 2414 2090 2418 2094
rect 2458 2090 2462 2094
rect 2508 2090 2512 2094
rect 2561 2090 2565 2094
rect 2590 2090 2594 2094
rect 2640 2090 2644 2094
rect 2693 2090 2697 2094
rect 2722 2090 2726 2094
rect 2772 2090 2776 2094
rect 2825 2090 2829 2094
rect 3248 2090 3252 2094
rect 3264 2090 3268 2096
rect 3298 2096 3302 2100
rect 3285 2090 3289 2094
rect 2296 2079 2300 2083
rect 2333 2077 2337 2081
rect 2353 2077 2357 2081
rect 2397 2077 2401 2081
rect 2481 2079 2485 2083
rect 1520 2060 1524 2064
rect 1536 2060 1540 2066
rect 1570 2066 1574 2070
rect 1557 2060 1561 2064
rect 1578 2060 1582 2064
rect 1594 2060 1598 2066
rect 1615 2060 1619 2064
rect 1631 2060 1635 2064
rect 1652 2060 1656 2064
rect 1668 2060 1672 2066
rect 1702 2066 1706 2070
rect 1689 2060 1693 2064
rect 1710 2060 1714 2064
rect 1726 2060 1730 2066
rect 1747 2060 1751 2064
rect 1763 2060 1767 2064
rect 1784 2060 1788 2064
rect 1800 2060 1804 2066
rect 1834 2066 1838 2070
rect 1821 2060 1825 2064
rect 1842 2060 1846 2064
rect 1858 2060 1862 2066
rect 1916 2070 1922 2074
rect 2452 2070 2456 2074
rect 2465 2073 2469 2079
rect 2502 2073 2506 2079
rect 2515 2075 2519 2079
rect 2539 2079 2543 2083
rect 2613 2079 2617 2083
rect 2523 2073 2527 2079
rect 2560 2073 2564 2079
rect 2576 2073 2580 2079
rect 2597 2073 2601 2079
rect 2634 2073 2638 2079
rect 2647 2075 2651 2079
rect 2671 2079 2675 2083
rect 2745 2079 2749 2083
rect 2655 2073 2659 2079
rect 2692 2073 2696 2079
rect 2708 2073 2712 2079
rect 2729 2073 2733 2079
rect 2766 2073 2770 2079
rect 2779 2075 2783 2079
rect 2803 2079 2807 2083
rect 2787 2073 2791 2079
rect 2824 2073 2828 2079
rect 2840 2075 2844 2079
rect 3306 2090 3310 2094
rect 3322 2090 3326 2096
rect 3343 2090 3347 2094
rect 3359 2090 3363 2094
rect 3241 2079 3245 2083
rect 3278 2077 3282 2081
rect 3298 2077 3302 2081
rect 3342 2077 3346 2081
rect 1879 2060 1883 2064
rect 1895 2060 1899 2064
rect 1952 2063 1958 2067
rect 2296 2063 2300 2067
rect 2347 2063 2351 2067
rect 2397 2063 2401 2067
rect 2465 2060 2469 2064
rect 2481 2060 2485 2066
rect 2515 2066 2519 2070
rect 2502 2060 2506 2064
rect 1513 2049 1517 2053
rect 1550 2047 1554 2051
rect 1570 2047 1574 2051
rect 1614 2047 1618 2051
rect 1645 2049 1649 2053
rect 1682 2047 1686 2051
rect 1702 2047 1706 2051
rect 1746 2047 1750 2051
rect 1777 2049 1781 2053
rect 1814 2047 1818 2051
rect 1834 2047 1838 2051
rect 1878 2047 1882 2051
rect 2289 2055 2293 2059
rect 2414 2056 2418 2060
rect 2523 2060 2527 2064
rect 2539 2060 2543 2066
rect 2560 2060 2564 2064
rect 2576 2060 2580 2064
rect 2597 2060 2601 2064
rect 2613 2060 2617 2066
rect 2647 2066 2651 2070
rect 2634 2060 2638 2064
rect 2655 2060 2659 2064
rect 2671 2060 2675 2066
rect 2692 2060 2696 2064
rect 2708 2060 2712 2064
rect 2729 2060 2733 2064
rect 2745 2060 2749 2066
rect 2779 2066 2783 2070
rect 2766 2060 2770 2064
rect 2787 2060 2791 2064
rect 2803 2060 2807 2066
rect 2861 2070 2867 2074
rect 2824 2060 2828 2064
rect 2840 2060 2844 2064
rect 2897 2063 2903 2067
rect 3241 2063 3245 2067
rect 3292 2063 3296 2067
rect 3342 2063 3346 2067
rect 1964 2048 1970 2052
rect 2296 2048 2300 2052
rect 2332 2048 2336 2052
rect 2399 2048 2403 2052
rect 1916 2040 1922 2044
rect 2282 2041 2286 2045
rect 2458 2049 2462 2053
rect 2495 2047 2499 2051
rect 2515 2047 2519 2051
rect 2559 2047 2563 2051
rect 2590 2049 2594 2053
rect 2627 2047 2631 2051
rect 2647 2047 2651 2051
rect 2691 2047 2695 2051
rect 2722 2049 2726 2053
rect 2759 2047 2763 2051
rect 2779 2047 2783 2051
rect 2823 2047 2827 2051
rect 3234 2055 3238 2059
rect 3359 2056 3363 2060
rect 2909 2048 2915 2052
rect 3241 2048 3245 2052
rect 3277 2048 3281 2052
rect 3344 2048 3348 2052
rect 1513 2033 1517 2037
rect 1564 2033 1568 2037
rect 1614 2033 1618 2037
rect 1645 2033 1649 2037
rect 1696 2033 1700 2037
rect 1746 2033 1750 2037
rect 1777 2033 1781 2037
rect 1828 2033 1832 2037
rect 1878 2033 1882 2037
rect 1952 2033 1958 2037
rect 2296 2034 2300 2038
rect 2346 2034 2350 2038
rect 2399 2034 2403 2038
rect 2861 2040 2867 2044
rect 3227 2041 3231 2045
rect 2458 2033 2462 2037
rect 2509 2033 2513 2037
rect 2559 2033 2563 2037
rect 2590 2033 2594 2037
rect 2641 2033 2645 2037
rect 2691 2033 2695 2037
rect 2722 2033 2726 2037
rect 2773 2033 2777 2037
rect 2823 2033 2827 2037
rect 2897 2033 2903 2037
rect 3241 2034 3245 2038
rect 3291 2034 3295 2038
rect 3344 2034 3348 2038
rect 1506 2026 1510 2030
rect 1895 2026 1899 2030
rect 2319 2023 2323 2027
rect 1513 2018 1517 2022
rect 1549 2018 1553 2022
rect 1616 2018 1620 2022
rect 1645 2018 1649 2022
rect 1681 2018 1685 2022
rect 1748 2018 1752 2022
rect 1777 2018 1781 2022
rect 1813 2018 1817 2022
rect 1880 2018 1884 2022
rect 1964 2018 1970 2022
rect 1904 2011 1910 2015
rect 2290 2014 2294 2018
rect 2303 2017 2307 2023
rect 2340 2017 2344 2023
rect 2353 2019 2357 2023
rect 2377 2023 2381 2027
rect 2451 2026 2455 2030
rect 2840 2026 2844 2030
rect 3264 2023 3268 2027
rect 2361 2017 2365 2023
rect 2398 2017 2402 2023
rect 2414 2019 2418 2023
rect 2436 2017 2440 2021
rect 2458 2018 2462 2022
rect 2494 2018 2498 2022
rect 2561 2018 2565 2022
rect 2590 2018 2594 2022
rect 2626 2018 2630 2022
rect 2693 2018 2697 2022
rect 2722 2018 2726 2022
rect 2758 2018 2762 2022
rect 2825 2018 2829 2022
rect 2909 2018 2915 2022
rect 1513 2004 1517 2008
rect 1563 2004 1567 2008
rect 1616 2004 1620 2008
rect 1645 2004 1649 2008
rect 1695 2004 1699 2008
rect 1748 2004 1752 2008
rect 1777 2004 1781 2008
rect 1827 2004 1831 2008
rect 1880 2004 1884 2008
rect 2303 2004 2307 2008
rect 2319 2004 2323 2010
rect 2353 2010 2357 2014
rect 2340 2004 2344 2008
rect 1536 1993 1540 1997
rect 1507 1984 1511 1988
rect 1520 1987 1524 1993
rect 1557 1987 1561 1993
rect 1570 1989 1574 1993
rect 1594 1993 1598 1997
rect 1668 1993 1672 1997
rect 1578 1987 1582 1993
rect 1615 1987 1619 1993
rect 1631 1987 1635 1993
rect 1652 1987 1656 1993
rect 1689 1987 1693 1993
rect 1702 1989 1706 1993
rect 1726 1993 1730 1997
rect 1800 1993 1804 1997
rect 1710 1987 1714 1993
rect 1747 1987 1751 1993
rect 1763 1987 1767 1993
rect 1784 1987 1788 1993
rect 1821 1987 1825 1993
rect 1834 1989 1838 1993
rect 1858 1993 1862 1997
rect 1842 1987 1846 1993
rect 1879 1987 1883 1993
rect 1895 1989 1899 1993
rect 2361 2004 2365 2008
rect 2377 2004 2381 2010
rect 2398 2004 2402 2008
rect 2414 2004 2418 2013
rect 2849 2011 2855 2015
rect 3235 2014 3239 2018
rect 3248 2017 3252 2023
rect 3285 2017 3289 2023
rect 3298 2019 3302 2023
rect 3322 2023 3326 2027
rect 3306 2017 3310 2023
rect 3343 2017 3347 2023
rect 3359 2019 3363 2023
rect 3381 2017 3385 2021
rect 2436 2001 2440 2005
rect 2458 2004 2462 2008
rect 2508 2004 2512 2008
rect 2561 2004 2565 2008
rect 2590 2004 2594 2008
rect 2640 2004 2644 2008
rect 2693 2004 2697 2008
rect 2722 2004 2726 2008
rect 2772 2004 2776 2008
rect 2825 2004 2829 2008
rect 3248 2004 3252 2008
rect 3264 2004 3268 2010
rect 3298 2010 3302 2014
rect 3285 2004 3289 2008
rect 2296 1993 2300 1997
rect 2333 1991 2337 1995
rect 2353 1991 2357 1995
rect 2397 1991 2401 1995
rect 2481 1993 2485 1997
rect 1520 1974 1524 1978
rect 1536 1974 1540 1980
rect 1570 1980 1574 1984
rect 1557 1974 1561 1978
rect 1578 1974 1582 1978
rect 1594 1974 1598 1980
rect 1615 1974 1619 1978
rect 1631 1974 1635 1978
rect 1652 1974 1656 1978
rect 1668 1974 1672 1980
rect 1702 1980 1706 1984
rect 1689 1974 1693 1978
rect 1710 1974 1714 1978
rect 1726 1974 1730 1980
rect 1747 1974 1751 1978
rect 1763 1974 1767 1978
rect 1784 1974 1788 1978
rect 1800 1974 1804 1980
rect 1834 1980 1838 1984
rect 1821 1974 1825 1978
rect 1842 1974 1846 1978
rect 1858 1974 1862 1980
rect 1916 1984 1922 1988
rect 2452 1984 2456 1988
rect 2465 1987 2469 1993
rect 2502 1987 2506 1993
rect 2515 1989 2519 1993
rect 2539 1993 2543 1997
rect 2613 1993 2617 1997
rect 2523 1987 2527 1993
rect 2560 1987 2564 1993
rect 2576 1987 2580 1993
rect 2597 1987 2601 1993
rect 2634 1987 2638 1993
rect 2647 1989 2651 1993
rect 2671 1993 2675 1997
rect 2745 1993 2749 1997
rect 2655 1987 2659 1993
rect 2692 1987 2696 1993
rect 2708 1987 2712 1993
rect 2729 1987 2733 1993
rect 2766 1987 2770 1993
rect 2779 1989 2783 1993
rect 2803 1993 2807 1997
rect 2787 1987 2791 1993
rect 2824 1987 2828 1993
rect 2840 1989 2844 1993
rect 3306 2004 3310 2008
rect 3322 2004 3326 2010
rect 3343 2004 3347 2008
rect 3359 2004 3363 2013
rect 3381 2001 3385 2005
rect 3241 1993 3245 1997
rect 3278 1991 3282 1995
rect 3298 1991 3302 1995
rect 3342 1991 3346 1995
rect 1879 1974 1883 1978
rect 1895 1974 1899 1978
rect 1952 1977 1958 1981
rect 2296 1977 2300 1981
rect 2347 1977 2351 1981
rect 2397 1977 2401 1981
rect 2465 1974 2469 1978
rect 2481 1974 2485 1980
rect 2515 1980 2519 1984
rect 2502 1974 2506 1978
rect 2523 1974 2527 1978
rect 2539 1974 2543 1980
rect 2560 1974 2564 1978
rect 2576 1974 2580 1978
rect 2597 1974 2601 1978
rect 2613 1974 2617 1980
rect 2647 1980 2651 1984
rect 2634 1974 2638 1978
rect 2655 1974 2659 1978
rect 2671 1974 2675 1980
rect 2692 1974 2696 1978
rect 2708 1974 2712 1978
rect 2729 1974 2733 1978
rect 2745 1974 2749 1980
rect 2779 1980 2783 1984
rect 2766 1974 2770 1978
rect 2787 1974 2791 1978
rect 2803 1974 2807 1980
rect 2861 1984 2867 1988
rect 2824 1974 2828 1978
rect 2840 1974 2844 1978
rect 2897 1977 2903 1981
rect 3241 1977 3245 1981
rect 3292 1977 3296 1981
rect 3342 1977 3346 1981
rect 1513 1963 1517 1967
rect 1550 1961 1554 1965
rect 1570 1961 1574 1965
rect 1614 1961 1618 1965
rect 1645 1963 1649 1967
rect 1682 1961 1686 1965
rect 1702 1961 1706 1965
rect 1746 1961 1750 1965
rect 1777 1963 1781 1967
rect 1814 1961 1818 1965
rect 1834 1961 1838 1965
rect 1878 1961 1882 1965
rect 2458 1963 2462 1967
rect 2495 1961 2499 1965
rect 2515 1961 2519 1965
rect 2559 1961 2563 1965
rect 2590 1963 2594 1967
rect 2627 1961 2631 1965
rect 2647 1961 2651 1965
rect 2691 1961 2695 1965
rect 2722 1963 2726 1967
rect 2759 1961 2763 1965
rect 2779 1961 2783 1965
rect 2823 1961 2827 1965
rect 1916 1954 1922 1958
rect 2861 1954 2867 1958
rect 1513 1947 1517 1951
rect 1564 1947 1568 1951
rect 1614 1947 1618 1951
rect 1645 1947 1649 1951
rect 1696 1947 1700 1951
rect 1746 1947 1750 1951
rect 1777 1947 1781 1951
rect 1828 1947 1832 1951
rect 1878 1947 1882 1951
rect 1952 1947 1958 1951
rect 2458 1947 2462 1951
rect 2509 1947 2513 1951
rect 2559 1947 2563 1951
rect 2590 1947 2594 1951
rect 2641 1947 2645 1951
rect 2691 1947 2695 1951
rect 2722 1947 2726 1951
rect 2773 1947 2777 1951
rect 2823 1947 2827 1951
rect 2897 1947 2903 1951
rect 1506 1940 1510 1944
rect 1895 1940 1899 1944
rect 2451 1940 2455 1944
rect 2840 1940 2844 1944
rect 1631 1933 1635 1937
rect 1739 1933 1743 1937
rect 1763 1933 1767 1937
rect 2576 1933 2580 1937
rect 2684 1933 2688 1937
rect 2708 1933 2712 1937
rect 1755 1926 1759 1930
rect 1739 1922 1743 1926
rect 1771 1922 1775 1926
rect 2700 1926 2704 1930
rect 2684 1922 2688 1926
rect 2716 1922 2720 1926
rect 1739 1915 1743 1919
rect 1771 1915 1775 1919
rect 2436 1915 2440 1919
rect 2684 1915 2688 1919
rect 2716 1915 2720 1919
rect 3381 1915 3385 1919
rect 1755 1908 1759 1912
rect 1895 1908 1899 1912
rect 2700 1908 2704 1912
rect 2840 1908 2844 1912
rect 1895 1900 1899 1904
rect 2840 1900 2844 1904
rect 1739 1896 1743 1900
rect 1771 1896 1775 1900
rect 1755 1892 1759 1896
rect 2684 1896 2688 1900
rect 2716 1896 2720 1900
rect 2700 1892 2704 1896
rect 1631 1885 1635 1889
rect 1739 1885 1743 1889
rect 1763 1885 1767 1889
rect 2576 1885 2580 1889
rect 2684 1885 2688 1889
rect 2708 1885 2712 1889
rect 1513 1878 1517 1882
rect 1549 1878 1553 1882
rect 1616 1878 1620 1882
rect 1645 1878 1649 1882
rect 1681 1878 1685 1882
rect 1748 1878 1752 1882
rect 1777 1878 1781 1882
rect 1813 1878 1817 1882
rect 1880 1878 1884 1882
rect 1964 1878 1970 1882
rect 2458 1878 2462 1882
rect 2494 1878 2498 1882
rect 2561 1878 2565 1882
rect 2590 1878 2594 1882
rect 2626 1878 2630 1882
rect 2693 1878 2697 1882
rect 2722 1878 2726 1882
rect 2758 1878 2762 1882
rect 2825 1878 2829 1882
rect 2909 1878 2915 1882
rect 1904 1871 1910 1875
rect 2849 1871 2855 1875
rect 1513 1864 1517 1868
rect 1563 1864 1567 1868
rect 1616 1864 1620 1868
rect 1645 1864 1649 1868
rect 1695 1864 1699 1868
rect 1748 1864 1752 1868
rect 1777 1864 1781 1868
rect 1827 1864 1831 1868
rect 1880 1864 1884 1868
rect 2458 1864 2462 1868
rect 2508 1864 2512 1868
rect 2561 1864 2565 1868
rect 2590 1864 2594 1868
rect 2640 1864 2644 1868
rect 2693 1864 2697 1868
rect 2722 1864 2726 1868
rect 2772 1864 2776 1868
rect 2825 1864 2829 1868
rect 1536 1853 1540 1857
rect 1507 1844 1511 1848
rect 1520 1847 1524 1853
rect 1557 1847 1561 1853
rect 1570 1849 1574 1853
rect 1594 1853 1598 1857
rect 1668 1853 1672 1857
rect 1578 1847 1582 1853
rect 1615 1847 1619 1853
rect 1631 1847 1635 1853
rect 1652 1847 1656 1853
rect 1689 1847 1693 1853
rect 1702 1849 1706 1853
rect 1726 1853 1730 1857
rect 1800 1853 1804 1857
rect 1710 1847 1714 1853
rect 1747 1847 1751 1853
rect 1763 1847 1767 1853
rect 1784 1847 1788 1853
rect 1821 1847 1825 1853
rect 1834 1849 1838 1853
rect 1858 1853 1862 1857
rect 2481 1853 2485 1857
rect 1842 1847 1846 1853
rect 1879 1847 1883 1853
rect 1895 1849 1899 1853
rect 1520 1834 1524 1838
rect 1536 1834 1540 1840
rect 1570 1840 1574 1844
rect 1557 1834 1561 1838
rect 1578 1834 1582 1838
rect 1594 1834 1598 1840
rect 1615 1834 1619 1838
rect 1631 1834 1635 1838
rect 1652 1834 1656 1838
rect 1668 1834 1672 1840
rect 1702 1840 1706 1844
rect 1689 1834 1693 1838
rect 1710 1834 1714 1838
rect 1726 1834 1730 1840
rect 1747 1834 1751 1838
rect 1763 1834 1767 1838
rect 1784 1834 1788 1838
rect 1800 1834 1804 1840
rect 1834 1840 1838 1844
rect 1821 1834 1825 1838
rect 1842 1834 1846 1838
rect 1858 1834 1862 1840
rect 2452 1844 2456 1848
rect 2465 1847 2469 1853
rect 2502 1847 2506 1853
rect 2515 1849 2519 1853
rect 2539 1853 2543 1857
rect 2613 1853 2617 1857
rect 2523 1847 2527 1853
rect 2560 1847 2564 1853
rect 2576 1847 2580 1853
rect 2597 1847 2601 1853
rect 2634 1847 2638 1853
rect 2647 1849 2651 1853
rect 2671 1853 2675 1857
rect 2745 1853 2749 1857
rect 2655 1847 2659 1853
rect 2692 1847 2696 1853
rect 2708 1847 2712 1853
rect 2729 1847 2733 1853
rect 2766 1847 2770 1853
rect 2779 1849 2783 1853
rect 2803 1853 2807 1857
rect 2787 1847 2791 1853
rect 2824 1847 2828 1853
rect 2840 1849 2844 1853
rect 1879 1834 1883 1838
rect 1895 1834 1899 1838
rect 2465 1834 2469 1838
rect 2481 1834 2485 1840
rect 2515 1840 2519 1844
rect 2502 1834 2506 1838
rect 2523 1834 2527 1838
rect 2539 1834 2543 1840
rect 2560 1834 2564 1838
rect 2576 1834 2580 1838
rect 2597 1834 2601 1838
rect 2613 1834 2617 1840
rect 2647 1840 2651 1844
rect 2634 1834 2638 1838
rect 2655 1834 2659 1838
rect 2671 1834 2675 1840
rect 2692 1834 2696 1838
rect 2708 1834 2712 1838
rect 2729 1834 2733 1838
rect 2745 1834 2749 1840
rect 2779 1840 2783 1844
rect 2766 1834 2770 1838
rect 2787 1834 2791 1838
rect 2803 1834 2807 1840
rect 2824 1834 2828 1838
rect 2840 1834 2844 1838
rect 1513 1823 1517 1827
rect 1550 1821 1554 1825
rect 1570 1821 1574 1825
rect 1614 1821 1618 1825
rect 1645 1823 1649 1827
rect 1682 1821 1686 1825
rect 1702 1821 1706 1825
rect 1746 1821 1750 1825
rect 1777 1823 1781 1827
rect 1814 1821 1818 1825
rect 1834 1821 1838 1825
rect 1878 1821 1882 1825
rect 2458 1823 2462 1827
rect 2495 1821 2499 1825
rect 2515 1821 2519 1825
rect 2559 1821 2563 1825
rect 2590 1823 2594 1827
rect 2627 1821 2631 1825
rect 2647 1821 2651 1825
rect 2691 1821 2695 1825
rect 2722 1823 2726 1827
rect 2759 1821 2763 1825
rect 2779 1821 2783 1825
rect 2823 1821 2827 1825
rect 1916 1814 1922 1818
rect 2861 1814 2867 1818
rect 1513 1807 1517 1811
rect 1564 1807 1568 1811
rect 1614 1807 1618 1811
rect 1645 1807 1649 1811
rect 1696 1807 1700 1811
rect 1746 1807 1750 1811
rect 1777 1807 1781 1811
rect 1828 1807 1832 1811
rect 1878 1807 1882 1811
rect 1952 1807 1958 1811
rect 2458 1807 2462 1811
rect 2509 1807 2513 1811
rect 2559 1807 2563 1811
rect 2590 1807 2594 1811
rect 2641 1807 2645 1811
rect 2691 1807 2695 1811
rect 2722 1807 2726 1811
rect 2773 1807 2777 1811
rect 2823 1807 2827 1811
rect 2897 1807 2903 1811
<< metal2 >>
rect 2080 4448 2088 4450
rect 2080 4443 2081 4448
rect 2086 4443 2088 4448
rect 2080 4330 2088 4443
rect 2080 4323 2093 4330
rect 2087 4300 2093 4323
rect 2171 4326 2172 4330
rect 2171 4300 2175 4326
rect 2027 3966 2040 4300
rect 1897 3819 1901 3962
rect 2336 3955 2349 4300
rect 2645 4196 2658 4312
rect 2691 4276 2694 4298
rect 2990 4294 2994 4299
rect 2691 4273 2736 4276
rect 2691 4263 2694 4273
rect 2669 4259 2690 4263
rect 2709 4260 2729 4263
rect 2645 4182 2660 4196
rect 2645 4178 2656 4182
rect 2656 4052 2660 4178
rect 2669 4133 2672 4259
rect 2691 4254 2694 4259
rect 2691 4251 2713 4254
rect 2726 4241 2729 4260
rect 2726 4161 2729 4237
rect 2737 4197 2740 4273
rect 2744 4181 2748 4251
rect 2691 4143 2736 4146
rect 2691 4133 2694 4143
rect 2709 4130 2729 4133
rect 2669 4124 2672 4129
rect 2669 4121 2713 4124
rect 2726 4111 2729 4130
rect 2656 4048 2658 4052
rect 2726 4031 2729 4107
rect 2737 4067 2740 4143
rect 2744 4051 2748 4121
rect 2866 4102 2903 4106
rect 2818 4064 2822 4101
rect 2818 4059 2891 4064
rect 1928 3925 1934 3947
rect 1616 3239 1620 3815
rect 1630 3647 1633 3696
rect 1630 3603 1633 3643
rect 1638 3640 1642 3807
rect 1646 3720 1649 3730
rect 1653 3690 1656 3699
rect 1669 3692 1672 3705
rect 1682 3677 1685 3730
rect 1749 3720 1752 3730
rect 1689 3705 1693 3709
rect 1690 3690 1693 3699
rect 1645 3663 1648 3675
rect 1686 3673 1687 3677
rect 1696 3663 1699 3716
rect 1702 3696 1705 3701
rect 1711 3690 1714 3699
rect 1727 3692 1730 3705
rect 1748 3690 1751 3699
rect 1747 3663 1750 3673
rect 1630 3588 1633 3597
rect 1491 3127 1495 3235
rect 1514 3218 1517 3228
rect 1521 3188 1524 3197
rect 1537 3190 1540 3203
rect 1550 3175 1553 3228
rect 1617 3218 1620 3228
rect 1557 3203 1561 3207
rect 1558 3188 1561 3197
rect 1513 3161 1516 3173
rect 1554 3171 1555 3175
rect 1564 3161 1567 3214
rect 1570 3194 1573 3199
rect 1579 3188 1582 3197
rect 1595 3190 1598 3203
rect 1616 3188 1619 3197
rect 1632 3188 1635 3197
rect 1615 3161 1618 3171
rect 1507 3056 1510 3150
rect 1632 3147 1635 3184
rect 1638 3140 1642 3636
rect 1755 3649 1759 3783
rect 1904 3760 1910 3905
rect 1904 3727 1910 3756
rect 1764 3697 1767 3699
rect 1764 3690 1767 3693
rect 1764 3656 1767 3686
rect 1904 3683 1910 3723
rect 1645 3618 1648 3628
rect 1646 3588 1649 3597
rect 1667 3590 1670 3603
rect 1683 3588 1686 3597
rect 1692 3594 1695 3599
rect 1647 3561 1650 3571
rect 1698 3561 1701 3614
rect 1704 3603 1708 3607
rect 1704 3588 1707 3597
rect 1712 3575 1715 3628
rect 1748 3618 1751 3628
rect 1725 3590 1728 3603
rect 1741 3588 1744 3597
rect 1710 3571 1711 3575
rect 1749 3561 1752 3573
rect 1646 3218 1649 3228
rect 1653 3188 1656 3197
rect 1669 3190 1672 3203
rect 1682 3175 1685 3228
rect 1749 3218 1752 3228
rect 1689 3203 1693 3207
rect 1690 3188 1693 3197
rect 1645 3161 1648 3173
rect 1686 3171 1687 3175
rect 1696 3161 1699 3214
rect 1702 3194 1705 3199
rect 1711 3188 1714 3197
rect 1727 3190 1730 3203
rect 1748 3188 1751 3197
rect 1747 3161 1750 3171
rect 1622 3127 1626 3131
rect 1622 3108 1626 3123
rect 1638 3120 1642 3136
rect 1654 3135 1658 3140
rect 1654 3127 1658 3131
rect 1654 3108 1658 3123
rect 1638 3104 1642 3105
rect 1654 3100 1658 3104
rect 1514 3076 1517 3086
rect 1521 3046 1524 3055
rect 1537 3048 1540 3061
rect 1550 3033 1553 3086
rect 1617 3076 1620 3086
rect 1557 3061 1561 3065
rect 1558 3046 1561 3055
rect 1513 3019 1516 3031
rect 1554 3029 1555 3033
rect 1564 3019 1567 3072
rect 1632 3061 1635 3093
rect 1570 3052 1573 3057
rect 1579 3046 1582 3055
rect 1595 3048 1598 3061
rect 1616 3046 1619 3055
rect 1632 3046 1635 3055
rect 1615 3019 1618 3029
rect 1507 2970 1510 3008
rect 1514 2990 1517 3000
rect 1521 2960 1524 2969
rect 1537 2962 1540 2975
rect 1550 2947 1553 3000
rect 1617 2990 1620 3000
rect 1557 2975 1561 2979
rect 1558 2960 1561 2969
rect 1513 2933 1516 2945
rect 1554 2943 1555 2947
rect 1564 2933 1567 2986
rect 1570 2966 1573 2971
rect 1579 2960 1582 2969
rect 1595 2962 1598 2975
rect 1616 2960 1619 2969
rect 1632 2960 1635 2969
rect 1615 2933 1618 2943
rect 1507 2830 1510 2922
rect 1632 2919 1635 2956
rect 1514 2850 1517 2860
rect 1521 2820 1524 2829
rect 1537 2822 1540 2835
rect 1550 2807 1553 2860
rect 1617 2850 1620 2860
rect 1557 2835 1561 2839
rect 1558 2820 1561 2829
rect 1513 2793 1516 2805
rect 1554 2803 1555 2807
rect 1564 2793 1567 2846
rect 1632 2835 1635 2867
rect 1570 2826 1573 2831
rect 1579 2820 1582 2829
rect 1595 2822 1598 2835
rect 1616 2820 1619 2829
rect 1632 2820 1635 2829
rect 1615 2793 1618 2803
rect 1630 2665 1633 2714
rect 1630 2621 1633 2661
rect 1638 2658 1642 3100
rect 1646 3076 1649 3086
rect 1653 3046 1656 3055
rect 1669 3048 1672 3061
rect 1682 3033 1685 3086
rect 1749 3076 1752 3086
rect 1689 3061 1693 3065
rect 1690 3046 1693 3055
rect 1645 3019 1648 3031
rect 1686 3029 1687 3033
rect 1696 3019 1699 3072
rect 1702 3052 1705 3057
rect 1711 3046 1714 3055
rect 1727 3048 1730 3061
rect 1748 3046 1751 3055
rect 1747 3019 1750 3029
rect 1646 2990 1649 3000
rect 1653 2960 1656 2969
rect 1669 2962 1672 2975
rect 1682 2947 1685 3000
rect 1749 2990 1752 3000
rect 1689 2975 1693 2979
rect 1690 2960 1693 2969
rect 1645 2933 1648 2945
rect 1686 2943 1687 2947
rect 1696 2933 1699 2986
rect 1702 2966 1705 2971
rect 1711 2960 1714 2969
rect 1727 2962 1730 2975
rect 1748 2960 1751 2969
rect 1747 2933 1750 2943
rect 1755 2912 1759 3645
rect 1779 3640 1783 3645
rect 1904 3625 1910 3679
rect 1904 3551 1910 3621
rect 1904 3419 1910 3547
rect 1904 3287 1910 3415
rect 1778 3218 1781 3228
rect 1764 3188 1767 3197
rect 1785 3188 1788 3197
rect 1801 3190 1804 3203
rect 1764 3147 1767 3184
rect 1814 3175 1817 3228
rect 1881 3218 1884 3228
rect 1904 3225 1910 3283
rect 1821 3203 1825 3207
rect 1822 3188 1825 3197
rect 1777 3161 1780 3173
rect 1818 3171 1819 3175
rect 1828 3161 1831 3214
rect 1834 3194 1837 3199
rect 1843 3188 1846 3197
rect 1859 3190 1862 3203
rect 1880 3188 1883 3197
rect 1896 3188 1899 3199
rect 1879 3161 1882 3171
rect 1896 3154 1899 3184
rect 1896 3120 1899 3150
rect 1904 3155 1910 3221
rect 1904 3113 1910 3151
rect 1764 3061 1767 3093
rect 1778 3076 1781 3086
rect 1764 3046 1767 3055
rect 1785 3046 1788 3055
rect 1801 3048 1804 3061
rect 1814 3033 1817 3086
rect 1881 3076 1884 3086
rect 1821 3061 1825 3065
rect 1822 3046 1825 3055
rect 1777 3019 1780 3031
rect 1818 3029 1819 3033
rect 1828 3019 1831 3072
rect 1896 3061 1899 3108
rect 1834 3052 1837 3057
rect 1843 3046 1846 3055
rect 1859 3048 1862 3061
rect 1880 3046 1883 3055
rect 1896 3046 1899 3057
rect 1879 3019 1882 3029
rect 1896 3012 1899 3042
rect 1904 3083 1910 3109
rect 1778 2990 1781 3000
rect 1764 2960 1767 2969
rect 1785 2960 1788 2969
rect 1801 2962 1804 2975
rect 1764 2919 1767 2956
rect 1814 2947 1817 3000
rect 1881 2990 1884 3000
rect 1904 2997 1910 3079
rect 1821 2975 1825 2979
rect 1822 2960 1825 2969
rect 1777 2933 1780 2945
rect 1818 2943 1819 2947
rect 1828 2933 1831 2986
rect 1834 2966 1837 2971
rect 1843 2960 1846 2969
rect 1859 2962 1862 2975
rect 1880 2960 1883 2969
rect 1896 2960 1899 2971
rect 1879 2933 1882 2943
rect 1896 2926 1899 2956
rect 1739 2901 1743 2904
rect 1739 2882 1743 2897
rect 1755 2894 1759 2908
rect 1771 2908 1775 2912
rect 1771 2901 1775 2904
rect 1771 2882 1775 2897
rect 1896 2894 1899 2922
rect 1755 2878 1759 2879
rect 1771 2874 1775 2878
rect 1646 2850 1649 2860
rect 1653 2820 1656 2829
rect 1669 2822 1672 2835
rect 1682 2807 1685 2860
rect 1749 2850 1752 2860
rect 1689 2835 1693 2839
rect 1690 2820 1693 2829
rect 1645 2793 1648 2805
rect 1686 2803 1687 2807
rect 1696 2793 1699 2846
rect 1702 2826 1705 2831
rect 1711 2820 1714 2829
rect 1727 2822 1730 2835
rect 1748 2820 1751 2829
rect 1747 2793 1750 2803
rect 1646 2738 1649 2748
rect 1653 2708 1656 2717
rect 1669 2710 1672 2723
rect 1682 2695 1685 2748
rect 1749 2738 1752 2748
rect 1689 2723 1693 2727
rect 1690 2708 1693 2717
rect 1645 2681 1648 2693
rect 1686 2691 1687 2695
rect 1696 2681 1699 2734
rect 1702 2714 1705 2719
rect 1711 2708 1714 2717
rect 1727 2710 1730 2723
rect 1748 2708 1751 2717
rect 1747 2681 1750 2691
rect 1630 2606 1633 2615
rect 1514 2236 1517 2246
rect 1521 2206 1524 2215
rect 1537 2208 1540 2221
rect 1550 2193 1553 2246
rect 1617 2236 1620 2246
rect 1557 2221 1561 2225
rect 1558 2206 1561 2215
rect 1513 2179 1516 2191
rect 1554 2189 1555 2193
rect 1564 2179 1567 2232
rect 1570 2212 1573 2217
rect 1579 2206 1582 2215
rect 1595 2208 1598 2221
rect 1616 2206 1619 2215
rect 1632 2206 1635 2215
rect 1615 2179 1618 2189
rect 1507 2074 1510 2168
rect 1632 2165 1635 2202
rect 1638 2158 1642 2654
rect 1755 2667 1759 2874
rect 1764 2835 1767 2867
rect 1778 2850 1781 2860
rect 1764 2820 1767 2829
rect 1785 2820 1788 2829
rect 1801 2822 1804 2835
rect 1814 2807 1817 2860
rect 1881 2850 1884 2860
rect 1821 2835 1825 2839
rect 1822 2820 1825 2829
rect 1777 2793 1780 2805
rect 1818 2803 1819 2807
rect 1828 2793 1831 2846
rect 1896 2835 1899 2882
rect 1834 2826 1837 2831
rect 1843 2820 1846 2829
rect 1859 2822 1862 2835
rect 1880 2820 1883 2829
rect 1896 2827 1899 2831
rect 1904 2857 1910 2993
rect 1896 2820 1899 2823
rect 1879 2793 1882 2803
rect 1904 2778 1910 2853
rect 1904 2745 1910 2774
rect 1764 2715 1767 2717
rect 1764 2708 1767 2711
rect 1764 2674 1767 2704
rect 1904 2701 1910 2741
rect 1645 2636 1648 2646
rect 1646 2606 1649 2615
rect 1667 2608 1670 2621
rect 1683 2606 1686 2615
rect 1692 2612 1695 2617
rect 1647 2579 1650 2589
rect 1698 2579 1701 2632
rect 1704 2621 1708 2625
rect 1704 2606 1707 2615
rect 1712 2593 1715 2646
rect 1748 2636 1751 2646
rect 1725 2608 1728 2621
rect 1741 2606 1744 2615
rect 1710 2589 1711 2593
rect 1749 2579 1752 2591
rect 1646 2236 1649 2246
rect 1653 2206 1656 2215
rect 1669 2208 1672 2221
rect 1682 2193 1685 2246
rect 1749 2236 1752 2246
rect 1689 2221 1693 2225
rect 1690 2206 1693 2215
rect 1645 2179 1648 2191
rect 1686 2189 1687 2193
rect 1696 2179 1699 2232
rect 1702 2212 1705 2217
rect 1711 2206 1714 2215
rect 1727 2208 1730 2221
rect 1748 2206 1751 2215
rect 1747 2179 1750 2189
rect 1622 2145 1626 2150
rect 1622 2126 1626 2141
rect 1638 2138 1642 2154
rect 1654 2154 1658 2158
rect 1654 2145 1658 2150
rect 1654 2126 1658 2141
rect 1638 2122 1642 2123
rect 1654 2118 1658 2122
rect 1514 2094 1517 2104
rect 1521 2064 1524 2073
rect 1537 2066 1540 2079
rect 1550 2051 1553 2104
rect 1617 2094 1620 2104
rect 1557 2079 1561 2083
rect 1558 2064 1561 2073
rect 1513 2037 1516 2049
rect 1554 2047 1555 2051
rect 1564 2037 1567 2090
rect 1632 2079 1635 2111
rect 1570 2070 1573 2075
rect 1579 2064 1582 2073
rect 1595 2066 1598 2079
rect 1616 2064 1619 2073
rect 1632 2064 1635 2073
rect 1615 2037 1618 2047
rect 1507 1988 1510 2026
rect 1514 2008 1517 2018
rect 1521 1978 1524 1987
rect 1537 1980 1540 1993
rect 1550 1965 1553 2018
rect 1617 2008 1620 2018
rect 1557 1993 1561 1997
rect 1558 1978 1561 1987
rect 1513 1951 1516 1963
rect 1554 1961 1555 1965
rect 1564 1951 1567 2004
rect 1570 1984 1573 1989
rect 1579 1978 1582 1987
rect 1595 1980 1598 1993
rect 1616 1978 1619 1987
rect 1632 1978 1635 1987
rect 1615 1951 1618 1961
rect 1507 1848 1510 1940
rect 1632 1937 1635 1974
rect 1514 1868 1517 1878
rect 1521 1838 1524 1847
rect 1537 1840 1540 1853
rect 1550 1825 1553 1878
rect 1617 1868 1620 1878
rect 1557 1853 1561 1857
rect 1558 1838 1561 1847
rect 1513 1811 1516 1823
rect 1554 1821 1555 1825
rect 1564 1811 1567 1864
rect 1632 1853 1635 1885
rect 1570 1844 1573 1849
rect 1579 1838 1582 1847
rect 1595 1840 1598 1853
rect 1616 1838 1619 1847
rect 1632 1838 1635 1847
rect 1615 1811 1618 1821
rect 1638 1797 1642 2118
rect 1646 2094 1649 2104
rect 1653 2064 1656 2073
rect 1669 2066 1672 2079
rect 1682 2051 1685 2104
rect 1749 2094 1752 2104
rect 1689 2079 1693 2083
rect 1690 2064 1693 2073
rect 1645 2037 1648 2049
rect 1686 2047 1687 2051
rect 1696 2037 1699 2090
rect 1702 2070 1705 2075
rect 1711 2064 1714 2073
rect 1727 2066 1730 2079
rect 1748 2064 1751 2073
rect 1747 2037 1750 2047
rect 1646 2008 1649 2018
rect 1653 1978 1656 1987
rect 1669 1980 1672 1993
rect 1682 1965 1685 2018
rect 1749 2008 1752 2018
rect 1689 1993 1693 1997
rect 1690 1978 1693 1987
rect 1645 1951 1648 1963
rect 1686 1961 1687 1965
rect 1696 1951 1699 2004
rect 1702 1984 1705 1989
rect 1711 1978 1714 1987
rect 1727 1980 1730 1993
rect 1748 1978 1751 1987
rect 1747 1951 1750 1961
rect 1755 1930 1759 2663
rect 1779 2658 1783 2663
rect 1904 2643 1910 2697
rect 1904 2569 1910 2639
rect 1904 2437 1910 2565
rect 1904 2305 1910 2433
rect 1778 2236 1781 2246
rect 1764 2206 1767 2215
rect 1785 2206 1788 2215
rect 1801 2208 1804 2221
rect 1764 2165 1767 2202
rect 1814 2193 1817 2246
rect 1881 2236 1884 2246
rect 1904 2243 1910 2301
rect 1821 2221 1825 2225
rect 1822 2206 1825 2215
rect 1777 2179 1780 2191
rect 1818 2189 1819 2193
rect 1828 2179 1831 2232
rect 1834 2212 1837 2217
rect 1843 2206 1846 2215
rect 1859 2208 1862 2221
rect 1880 2206 1883 2215
rect 1896 2206 1899 2217
rect 1879 2179 1882 2189
rect 1896 2172 1899 2202
rect 1896 2138 1899 2168
rect 1904 2173 1910 2239
rect 1904 2131 1910 2169
rect 1764 2079 1767 2111
rect 1778 2094 1781 2104
rect 1764 2064 1767 2073
rect 1785 2064 1788 2073
rect 1801 2066 1804 2079
rect 1814 2051 1817 2104
rect 1881 2094 1884 2104
rect 1821 2079 1825 2083
rect 1822 2064 1825 2073
rect 1777 2037 1780 2049
rect 1818 2047 1819 2051
rect 1828 2037 1831 2090
rect 1896 2079 1899 2126
rect 1834 2070 1837 2075
rect 1843 2064 1846 2073
rect 1859 2066 1862 2079
rect 1880 2064 1883 2073
rect 1896 2064 1899 2075
rect 1879 2037 1882 2047
rect 1896 2030 1899 2060
rect 1904 2101 1910 2127
rect 1778 2008 1781 2018
rect 1764 1978 1767 1987
rect 1785 1978 1788 1987
rect 1801 1980 1804 1993
rect 1764 1937 1767 1974
rect 1814 1965 1817 2018
rect 1881 2008 1884 2018
rect 1904 2015 1910 2097
rect 1821 1993 1825 1997
rect 1822 1978 1825 1987
rect 1777 1951 1780 1963
rect 1818 1961 1819 1965
rect 1828 1951 1831 2004
rect 1834 1984 1837 1989
rect 1843 1978 1846 1987
rect 1859 1980 1862 1993
rect 1880 1978 1883 1987
rect 1896 1978 1899 1989
rect 1879 1951 1882 1961
rect 1896 1944 1899 1974
rect 1739 1919 1743 1922
rect 1739 1900 1743 1915
rect 1755 1912 1759 1926
rect 1771 1926 1775 1930
rect 1771 1919 1775 1922
rect 1771 1900 1775 1915
rect 1896 1912 1899 1940
rect 1755 1896 1759 1897
rect 1771 1892 1775 1896
rect 1646 1868 1649 1878
rect 1653 1838 1656 1847
rect 1669 1840 1672 1853
rect 1682 1825 1685 1878
rect 1749 1868 1752 1878
rect 1689 1853 1693 1857
rect 1690 1838 1693 1847
rect 1645 1811 1648 1823
rect 1686 1821 1687 1825
rect 1696 1811 1699 1864
rect 1702 1844 1705 1849
rect 1711 1838 1714 1847
rect 1727 1840 1730 1853
rect 1748 1838 1751 1847
rect 1747 1811 1750 1821
rect 1755 1797 1759 1892
rect 1764 1853 1767 1885
rect 1778 1868 1781 1878
rect 1764 1838 1767 1847
rect 1785 1838 1788 1847
rect 1801 1840 1804 1853
rect 1814 1825 1817 1878
rect 1881 1868 1884 1878
rect 1821 1853 1825 1857
rect 1822 1838 1825 1847
rect 1777 1811 1780 1823
rect 1818 1821 1819 1825
rect 1828 1811 1831 1864
rect 1896 1853 1899 1900
rect 1834 1844 1837 1849
rect 1843 1838 1846 1847
rect 1859 1840 1862 1853
rect 1880 1838 1883 1847
rect 1896 1845 1899 1849
rect 1904 1875 1910 2011
rect 1896 1838 1899 1841
rect 1879 1811 1882 1821
rect 1904 1797 1910 1871
rect 1916 3703 1922 3912
rect 1916 3670 1922 3699
rect 1916 3617 1922 3666
rect 1916 3568 1922 3613
rect 1916 3485 1922 3564
rect 1916 3353 1922 3481
rect 1916 3221 1922 3349
rect 1916 3168 1922 3217
rect 1916 3056 1922 3164
rect 1916 3026 1922 3052
rect 1916 2970 1922 3022
rect 1916 2940 1922 2966
rect 1916 2800 1922 2936
rect 1916 2721 1922 2796
rect 1916 2688 1922 2717
rect 1916 2635 1922 2684
rect 1916 2586 1922 2631
rect 1916 2503 1922 2582
rect 1916 2371 1922 2499
rect 1916 2239 1922 2367
rect 1916 2186 1922 2235
rect 1916 2074 1922 2182
rect 1916 2044 1922 2070
rect 1916 1988 1922 2040
rect 1916 1958 1922 1984
rect 1916 1818 1922 1954
rect 1916 1797 1922 1814
rect 1928 3624 1934 3921
rect 1928 3610 1934 3620
rect 1928 3492 1934 3606
rect 1928 3478 1934 3488
rect 1928 3360 1934 3474
rect 1928 3346 1934 3356
rect 1928 3214 1934 3342
rect 1928 3140 1934 3210
rect 1928 2642 1934 3136
rect 1928 2628 1934 2638
rect 1928 2510 1934 2624
rect 1928 2496 1934 2506
rect 1928 2378 1934 2492
rect 1928 2364 1934 2374
rect 1928 2232 1934 2360
rect 1928 2158 1934 2228
rect 1928 1797 1934 2154
rect 1940 3932 1946 3947
rect 1940 3676 1946 3928
rect 1940 3544 1946 3672
rect 1940 3426 1946 3540
rect 1940 3412 1946 3422
rect 1940 3294 1946 3408
rect 1940 3280 1946 3290
rect 1940 3148 1946 3276
rect 1940 2694 1946 3144
rect 1940 2562 1946 2690
rect 1940 2444 1946 2558
rect 1940 2430 1946 2440
rect 1940 2312 1946 2426
rect 1940 2298 1946 2308
rect 1940 2166 1946 2294
rect 1940 1797 1946 2162
rect 1952 3939 1958 3947
rect 1952 3696 1958 3935
rect 1952 3663 1958 3692
rect 1952 3561 1958 3659
rect 1952 3162 1958 3557
rect 1952 3049 1958 3158
rect 1952 3019 1958 3045
rect 1952 2963 1958 3015
rect 1952 2933 1958 2959
rect 1952 2793 1958 2929
rect 1952 2714 1958 2789
rect 1952 2681 1958 2710
rect 1952 2579 1958 2677
rect 1952 2180 1958 2575
rect 1952 2067 1958 2176
rect 1952 2037 1958 2063
rect 1952 1981 1958 2033
rect 1952 1951 1958 1977
rect 1952 1811 1958 1947
rect 1952 1797 1958 1807
rect 1964 3767 1970 3943
rect 1964 3734 1970 3763
rect 1964 3632 1970 3730
rect 1964 3232 1970 3628
rect 1964 3120 1970 3228
rect 1964 3090 1970 3116
rect 1964 3034 1970 3086
rect 1964 3004 1970 3030
rect 1964 2864 1970 3000
rect 1964 2785 1970 2860
rect 1964 2752 1970 2781
rect 1964 2650 1970 2748
rect 1964 2250 1970 2646
rect 1964 2138 1970 2246
rect 1964 2108 1970 2134
rect 1964 2052 1970 2104
rect 1964 2022 1970 2048
rect 1964 1882 1970 2018
rect 1964 1797 1970 1878
rect 1976 3134 1982 3898
rect 1987 3811 1991 3951
rect 2861 3925 2867 3994
rect 2837 3800 2843 3906
rect 2849 3808 2855 3913
rect 2849 3800 2855 3804
rect 1998 3753 2001 3763
rect 1987 3733 1991 3734
rect 2005 3723 2008 3732
rect 2021 3725 2024 3738
rect 2034 3710 2037 3763
rect 2101 3753 2104 3763
rect 2130 3753 2133 3763
rect 2041 3738 2045 3742
rect 2042 3723 2045 3732
rect 1997 3696 2000 3708
rect 2038 3706 2039 3710
rect 2048 3696 2051 3749
rect 2054 3729 2057 3734
rect 2063 3723 2066 3732
rect 2079 3725 2082 3738
rect 2100 3723 2103 3732
rect 2116 3732 2119 3734
rect 2116 3729 2123 3732
rect 2116 3723 2119 3729
rect 2137 3723 2140 3732
rect 2153 3725 2156 3738
rect 2099 3696 2102 3706
rect 2116 3689 2119 3719
rect 2166 3710 2169 3763
rect 2233 3753 2236 3763
rect 2262 3753 2265 3763
rect 2173 3738 2177 3742
rect 2174 3723 2177 3732
rect 2129 3696 2132 3708
rect 2170 3706 2171 3710
rect 2180 3696 2183 3749
rect 2186 3729 2189 3734
rect 2195 3723 2198 3732
rect 2211 3725 2214 3738
rect 2232 3723 2235 3732
rect 2248 3732 2251 3734
rect 2248 3729 2255 3732
rect 2248 3723 2251 3729
rect 2269 3723 2272 3732
rect 2285 3725 2288 3738
rect 2231 3696 2234 3706
rect 2116 3686 2168 3689
rect 1996 3666 1999 3679
rect 2022 3669 2025 3672
rect 2029 3666 2032 3679
rect 2046 3666 2049 3679
rect 1996 3617 1999 3632
rect 2010 3624 2013 3628
rect 2028 3617 2031 3632
rect 2047 3617 2050 3632
rect 2053 3631 2056 3672
rect 2069 3624 2072 3665
rect 2075 3632 2078 3672
rect 2094 3624 2097 3665
rect 2103 3666 2106 3679
rect 2119 3666 2122 3679
rect 2140 3669 2143 3672
rect 2147 3666 2150 3679
rect 2165 3675 2168 3686
rect 2248 3683 2251 3719
rect 2298 3710 2301 3763
rect 2365 3753 2368 3763
rect 2394 3753 2397 3763
rect 2305 3738 2309 3742
rect 2306 3723 2309 3732
rect 2261 3696 2264 3708
rect 2302 3706 2303 3710
rect 2312 3696 2315 3749
rect 2318 3729 2321 3734
rect 2327 3723 2330 3732
rect 2343 3725 2346 3738
rect 2364 3723 2367 3732
rect 2380 3732 2383 3734
rect 2380 3729 2387 3732
rect 2380 3723 2383 3729
rect 2401 3723 2404 3732
rect 2417 3725 2420 3738
rect 2363 3696 2366 3706
rect 2380 3689 2383 3711
rect 2430 3710 2433 3763
rect 2497 3753 2500 3763
rect 2437 3738 2441 3742
rect 2438 3723 2441 3732
rect 2393 3696 2396 3708
rect 2434 3706 2435 3710
rect 2444 3696 2447 3749
rect 2450 3729 2453 3734
rect 2459 3723 2462 3732
rect 2475 3725 2478 3738
rect 2496 3723 2499 3732
rect 2512 3732 2515 3734
rect 2512 3729 2516 3732
rect 2512 3723 2515 3729
rect 2512 3715 2515 3719
rect 2495 3696 2498 3706
rect 2246 3678 2251 3683
rect 2308 3685 2383 3689
rect 2165 3672 2210 3675
rect 2165 3662 2168 3672
rect 2183 3659 2203 3662
rect 2200 3640 2203 3659
rect 2103 3617 2106 3632
rect 2118 3617 2121 3632
rect 2125 3624 2129 3627
rect 2146 3617 2149 3632
rect 1996 3598 1999 3613
rect 2010 3602 2013 3606
rect 2028 3598 2031 3613
rect 2047 3598 2050 3613
rect 1996 3551 1999 3564
rect 2022 3558 2025 3561
rect 1996 3534 1999 3547
rect 2006 3544 2010 3554
rect 2029 3551 2032 3564
rect 2046 3551 2049 3564
rect 2053 3558 2056 3599
rect 2069 3565 2072 3606
rect 2075 3558 2078 3598
rect 2094 3565 2097 3606
rect 2103 3598 2106 3613
rect 2118 3598 2121 3613
rect 2125 3603 2129 3606
rect 2146 3598 2149 3613
rect 2103 3551 2106 3564
rect 2022 3537 2025 3540
rect 2029 3534 2032 3547
rect 2046 3534 2049 3547
rect 1996 3485 1999 3500
rect 2010 3492 2013 3496
rect 2028 3485 2031 3500
rect 2047 3485 2050 3500
rect 2053 3499 2056 3540
rect 2069 3492 2072 3533
rect 2075 3500 2078 3540
rect 2094 3492 2097 3533
rect 2103 3534 2106 3547
rect 2119 3551 2122 3564
rect 2140 3558 2143 3561
rect 2147 3551 2150 3564
rect 2200 3564 2203 3636
rect 2211 3600 2214 3672
rect 2246 3675 2249 3678
rect 2246 3672 2291 3675
rect 2246 3662 2249 3672
rect 2119 3534 2122 3547
rect 2140 3537 2143 3540
rect 2147 3534 2150 3547
rect 2200 3530 2203 3560
rect 2211 3544 2214 3596
rect 2218 3584 2222 3650
rect 2206 3540 2210 3543
rect 2199 3527 2203 3530
rect 2200 3508 2203 3527
rect 2103 3485 2106 3500
rect 2118 3485 2121 3500
rect 2125 3492 2129 3495
rect 2146 3485 2149 3500
rect 1996 3466 1999 3481
rect 2010 3470 2013 3474
rect 2028 3466 2031 3481
rect 2047 3466 2050 3481
rect 1996 3419 1999 3432
rect 2022 3426 2025 3429
rect 1996 3402 1999 3415
rect 2029 3419 2032 3432
rect 2046 3419 2049 3432
rect 2053 3426 2056 3467
rect 2069 3433 2072 3474
rect 2075 3426 2078 3466
rect 2094 3433 2097 3474
rect 2103 3466 2106 3481
rect 2118 3466 2121 3481
rect 2125 3471 2129 3474
rect 2146 3466 2149 3481
rect 2103 3419 2106 3432
rect 2022 3405 2025 3408
rect 2029 3402 2032 3415
rect 2046 3402 2049 3415
rect 1996 3353 1999 3368
rect 2010 3360 2013 3364
rect 2028 3353 2031 3368
rect 2047 3353 2050 3368
rect 2053 3367 2056 3408
rect 2069 3360 2072 3401
rect 2075 3368 2078 3408
rect 2094 3360 2097 3401
rect 2103 3402 2106 3415
rect 2119 3419 2122 3432
rect 2140 3426 2143 3429
rect 2147 3419 2150 3432
rect 2200 3433 2203 3504
rect 2211 3469 2214 3540
rect 2119 3402 2122 3415
rect 2140 3405 2143 3408
rect 2147 3402 2150 3415
rect 2200 3376 2203 3429
rect 2211 3412 2214 3465
rect 2218 3453 2222 3518
rect 2206 3408 2210 3411
rect 2249 3411 2252 3662
rect 2264 3659 2284 3662
rect 2281 3640 2284 3659
rect 2281 3564 2284 3636
rect 2292 3600 2295 3672
rect 2299 3584 2303 3650
rect 2308 3551 2311 3685
rect 2512 3682 2515 3711
rect 2336 3679 2443 3682
rect 2270 3547 2311 3551
rect 2270 3543 2273 3547
rect 2270 3540 2315 3543
rect 2270 3530 2273 3540
rect 2288 3527 2308 3530
rect 2270 3525 2273 3526
rect 2305 3508 2308 3527
rect 2305 3433 2308 3504
rect 2316 3469 2319 3540
rect 2323 3453 2327 3518
rect 2103 3353 2106 3368
rect 2118 3353 2121 3368
rect 2125 3360 2129 3363
rect 2146 3353 2149 3368
rect 1996 3334 1999 3349
rect 2010 3338 2013 3342
rect 2028 3334 2031 3349
rect 2047 3334 2050 3349
rect 1996 3287 1999 3300
rect 2022 3294 2025 3297
rect 1996 3270 1999 3283
rect 2029 3287 2032 3300
rect 2046 3287 2049 3300
rect 2053 3294 2056 3335
rect 2069 3301 2072 3342
rect 2075 3294 2078 3334
rect 2094 3301 2097 3342
rect 2103 3334 2106 3349
rect 2118 3334 2121 3349
rect 2125 3339 2129 3342
rect 2146 3334 2149 3349
rect 2103 3287 2106 3300
rect 2022 3273 2025 3276
rect 2029 3270 2032 3283
rect 2046 3270 2049 3283
rect 1996 3221 1999 3236
rect 2010 3228 2013 3232
rect 1996 3202 1999 3217
rect 2019 3214 2023 3224
rect 2028 3221 2031 3236
rect 2047 3221 2050 3236
rect 2053 3235 2056 3276
rect 2069 3228 2072 3269
rect 2075 3236 2078 3276
rect 2094 3228 2097 3269
rect 2103 3270 2106 3283
rect 2119 3287 2122 3300
rect 2140 3294 2143 3297
rect 2147 3287 2150 3300
rect 2200 3298 2203 3372
rect 2211 3334 2214 3408
rect 2246 3408 2291 3411
rect 2246 3398 2249 3408
rect 2264 3395 2284 3398
rect 2119 3270 2122 3283
rect 2140 3273 2143 3276
rect 2147 3270 2150 3283
rect 2200 3244 2203 3294
rect 2211 3280 2214 3330
rect 2218 3318 2222 3386
rect 2281 3376 2284 3395
rect 2281 3298 2284 3372
rect 2292 3334 2295 3408
rect 2336 3411 2339 3679
rect 2447 3679 2515 3682
rect 2575 3647 2578 3696
rect 2575 3603 2578 3643
rect 2583 3640 2587 3783
rect 2591 3720 2594 3730
rect 2598 3690 2601 3699
rect 2614 3692 2617 3705
rect 2627 3677 2630 3730
rect 2694 3720 2697 3730
rect 2634 3705 2638 3709
rect 2635 3690 2638 3699
rect 2590 3663 2593 3675
rect 2631 3673 2632 3677
rect 2641 3663 2644 3716
rect 2647 3696 2650 3701
rect 2656 3690 2659 3699
rect 2672 3692 2675 3705
rect 2693 3690 2696 3699
rect 2692 3663 2695 3673
rect 2575 3588 2578 3597
rect 2336 3408 2381 3411
rect 2336 3398 2339 3408
rect 2354 3395 2374 3398
rect 2299 3318 2303 3386
rect 2371 3376 2374 3395
rect 2371 3298 2374 3372
rect 2382 3334 2385 3408
rect 2389 3318 2393 3386
rect 2206 3276 2210 3279
rect 2103 3221 2106 3236
rect 2118 3221 2121 3236
rect 2125 3228 2129 3231
rect 2146 3221 2149 3236
rect 2010 3206 2013 3210
rect 2028 3202 2031 3217
rect 2047 3202 2050 3217
rect 1996 3155 1999 3168
rect 2022 3162 2025 3165
rect 2004 3148 2008 3158
rect 2029 3155 2032 3168
rect 2046 3155 2049 3168
rect 2053 3162 2056 3203
rect 2069 3169 2072 3210
rect 2075 3162 2078 3202
rect 2094 3169 2097 3210
rect 2103 3202 2106 3217
rect 2118 3202 2121 3217
rect 2125 3207 2129 3210
rect 2146 3202 2149 3217
rect 2103 3155 2106 3168
rect 2119 3155 2122 3168
rect 2140 3162 2143 3165
rect 2147 3155 2150 3168
rect 2200 3162 2203 3240
rect 2211 3198 2214 3276
rect 2218 3182 2222 3254
rect 2230 3155 2234 3168
rect 2239 3148 2242 3158
rect 2249 3141 2252 3210
rect 2271 3206 2274 3210
rect 2289 3202 2292 3217
rect 2308 3202 2311 3217
rect 2256 3155 2260 3168
rect 2283 3162 2286 3165
rect 2290 3155 2293 3168
rect 2307 3155 2310 3168
rect 2314 3162 2317 3203
rect 2330 3169 2333 3210
rect 2336 3162 2339 3202
rect 2355 3169 2358 3210
rect 2364 3202 2367 3217
rect 2379 3202 2382 3217
rect 2386 3207 2390 3210
rect 2407 3202 2410 3217
rect 2364 3155 2367 3168
rect 2380 3155 2383 3168
rect 2401 3162 2404 3165
rect 2408 3155 2411 3168
rect 2424 3149 2428 3385
rect 2459 3218 2462 3228
rect 2466 3188 2469 3197
rect 2482 3190 2485 3203
rect 2495 3175 2498 3228
rect 2562 3218 2565 3228
rect 2502 3203 2506 3207
rect 2503 3188 2506 3197
rect 2458 3161 2461 3173
rect 2499 3171 2500 3175
rect 2509 3161 2512 3214
rect 2515 3194 2518 3199
rect 2524 3188 2527 3197
rect 2540 3190 2543 3203
rect 2561 3188 2564 3197
rect 2577 3188 2580 3197
rect 2560 3161 2563 3171
rect 2417 3137 2418 3140
rect 1976 2152 1982 3130
rect 2282 3027 2286 3109
rect 2297 3106 2300 3116
rect 2304 3076 2307 3085
rect 2320 3078 2323 3091
rect 2333 3063 2336 3116
rect 2400 3106 2403 3116
rect 2340 3091 2344 3095
rect 2341 3076 2344 3085
rect 2296 3049 2299 3061
rect 2337 3059 2338 3063
rect 2347 3049 2350 3102
rect 2415 3091 2418 3137
rect 2353 3082 2356 3087
rect 2362 3076 2365 3085
rect 2378 3078 2381 3091
rect 2399 3076 2402 3085
rect 2415 3076 2418 3085
rect 2398 3049 2401 3059
rect 2415 3042 2418 3072
rect 2290 3000 2293 3037
rect 2297 3020 2300 3030
rect 2304 2990 2307 2999
rect 2320 2992 2323 3005
rect 2333 2977 2336 3030
rect 2400 3020 2403 3030
rect 2340 3005 2344 3009
rect 2341 2990 2344 2999
rect 2296 2963 2299 2975
rect 2337 2973 2338 2977
rect 2347 2963 2350 3016
rect 2353 2996 2356 3001
rect 2362 2990 2365 2999
rect 2378 2992 2381 3005
rect 2399 2990 2402 2999
rect 2415 3000 2418 3001
rect 2436 3003 2440 3145
rect 2452 3056 2455 3150
rect 2577 3147 2580 3184
rect 2583 3140 2587 3636
rect 2700 3649 2704 3783
rect 2849 3760 2855 3796
rect 2849 3727 2855 3756
rect 2709 3697 2712 3699
rect 2709 3690 2712 3693
rect 2709 3656 2712 3686
rect 2849 3683 2855 3723
rect 2590 3618 2593 3628
rect 2591 3588 2594 3597
rect 2612 3590 2615 3603
rect 2628 3588 2631 3597
rect 2637 3594 2640 3599
rect 2592 3561 2595 3571
rect 2643 3561 2646 3614
rect 2649 3603 2653 3607
rect 2649 3588 2652 3597
rect 2657 3575 2660 3628
rect 2693 3618 2696 3628
rect 2670 3590 2673 3603
rect 2686 3588 2689 3597
rect 2655 3571 2656 3575
rect 2694 3561 2697 3573
rect 2591 3218 2594 3228
rect 2598 3188 2601 3197
rect 2614 3190 2617 3203
rect 2627 3175 2630 3228
rect 2694 3218 2697 3228
rect 2634 3203 2638 3207
rect 2635 3188 2638 3197
rect 2590 3161 2593 3173
rect 2631 3171 2632 3175
rect 2641 3161 2644 3214
rect 2647 3194 2650 3199
rect 2656 3188 2659 3197
rect 2672 3190 2675 3203
rect 2693 3188 2696 3197
rect 2692 3161 2695 3171
rect 2567 3127 2571 3131
rect 2567 3108 2571 3123
rect 2583 3120 2587 3136
rect 2599 3135 2603 3140
rect 2599 3127 2603 3131
rect 2599 3108 2603 3123
rect 2583 3104 2587 3105
rect 2599 3100 2603 3104
rect 2459 3076 2462 3086
rect 2466 3046 2469 3055
rect 2482 3048 2485 3061
rect 2495 3033 2498 3086
rect 2562 3076 2565 3086
rect 2502 3061 2506 3065
rect 2503 3046 2506 3055
rect 2458 3019 2461 3031
rect 2499 3029 2500 3033
rect 2509 3019 2512 3072
rect 2577 3061 2580 3093
rect 2515 3052 2518 3057
rect 2524 3046 2527 3055
rect 2540 3048 2543 3061
rect 2561 3046 2564 3055
rect 2577 3046 2580 3055
rect 2560 3019 2563 3029
rect 2415 2995 2418 2996
rect 2398 2963 2401 2973
rect 2436 2901 2440 2983
rect 2452 2970 2455 3008
rect 2459 2990 2462 3000
rect 2466 2960 2469 2969
rect 2482 2962 2485 2975
rect 2495 2947 2498 3000
rect 2562 2990 2565 3000
rect 2502 2975 2506 2979
rect 2503 2960 2506 2969
rect 2458 2933 2461 2945
rect 2499 2943 2500 2947
rect 2509 2933 2512 2986
rect 2515 2966 2518 2971
rect 2524 2960 2527 2969
rect 2540 2962 2543 2975
rect 2561 2960 2564 2969
rect 2577 2960 2580 2969
rect 2560 2933 2563 2943
rect 2452 2830 2455 2922
rect 2577 2919 2580 2956
rect 2459 2850 2462 2860
rect 2466 2820 2469 2829
rect 2482 2822 2485 2835
rect 2495 2807 2498 2860
rect 2562 2850 2565 2860
rect 2502 2835 2506 2839
rect 2503 2820 2506 2829
rect 2458 2793 2461 2805
rect 2499 2803 2500 2807
rect 2509 2793 2512 2846
rect 2577 2835 2580 2867
rect 2515 2826 2518 2831
rect 2524 2820 2527 2829
rect 2540 2822 2543 2835
rect 2561 2820 2564 2829
rect 2577 2820 2580 2829
rect 2560 2793 2563 2803
rect 1998 2771 2001 2781
rect 2005 2741 2008 2750
rect 2021 2743 2024 2756
rect 2034 2728 2037 2781
rect 2101 2771 2104 2781
rect 2130 2771 2133 2781
rect 2041 2756 2045 2760
rect 2042 2741 2045 2750
rect 1997 2714 2000 2726
rect 2038 2724 2039 2728
rect 2048 2714 2051 2767
rect 2054 2747 2057 2752
rect 2063 2741 2066 2750
rect 2079 2743 2082 2756
rect 2100 2741 2103 2750
rect 2116 2750 2119 2752
rect 2116 2747 2123 2750
rect 2116 2741 2119 2747
rect 2137 2741 2140 2750
rect 2153 2743 2156 2756
rect 2099 2714 2102 2724
rect 2116 2707 2119 2737
rect 2166 2728 2169 2781
rect 2233 2771 2236 2781
rect 2262 2771 2265 2781
rect 2173 2756 2177 2760
rect 2174 2741 2177 2750
rect 2129 2714 2132 2726
rect 2170 2724 2171 2728
rect 2180 2714 2183 2767
rect 2186 2747 2189 2752
rect 2195 2741 2198 2750
rect 2211 2743 2214 2756
rect 2232 2741 2235 2750
rect 2248 2750 2251 2752
rect 2248 2747 2255 2750
rect 2248 2741 2251 2747
rect 2269 2741 2272 2750
rect 2285 2743 2288 2756
rect 2231 2714 2234 2724
rect 2116 2704 2168 2707
rect 1996 2684 1999 2697
rect 2022 2687 2025 2690
rect 2029 2684 2032 2697
rect 2046 2684 2049 2697
rect 1996 2635 1999 2650
rect 2010 2642 2013 2646
rect 2028 2635 2031 2650
rect 2047 2635 2050 2650
rect 2053 2649 2056 2690
rect 2069 2642 2072 2683
rect 2075 2650 2078 2690
rect 2094 2642 2097 2683
rect 2103 2684 2106 2697
rect 2119 2684 2122 2697
rect 2140 2687 2143 2690
rect 2147 2684 2150 2697
rect 2165 2693 2168 2704
rect 2248 2701 2251 2737
rect 2298 2728 2301 2781
rect 2365 2771 2368 2781
rect 2394 2771 2397 2781
rect 2305 2756 2309 2760
rect 2306 2741 2309 2750
rect 2261 2714 2264 2726
rect 2302 2724 2303 2728
rect 2312 2714 2315 2767
rect 2318 2747 2321 2752
rect 2327 2741 2330 2750
rect 2343 2743 2346 2756
rect 2364 2741 2367 2750
rect 2380 2750 2383 2752
rect 2380 2747 2387 2750
rect 2380 2741 2383 2747
rect 2401 2741 2404 2750
rect 2417 2743 2420 2756
rect 2363 2714 2366 2724
rect 2380 2707 2383 2729
rect 2430 2728 2433 2781
rect 2497 2771 2500 2781
rect 2437 2756 2441 2760
rect 2438 2741 2441 2750
rect 2393 2714 2396 2726
rect 2434 2724 2435 2728
rect 2444 2714 2447 2767
rect 2450 2747 2453 2752
rect 2459 2741 2462 2750
rect 2475 2743 2478 2756
rect 2496 2741 2499 2750
rect 2512 2750 2515 2752
rect 2512 2747 2516 2750
rect 2512 2741 2515 2747
rect 2512 2733 2515 2737
rect 2495 2714 2498 2724
rect 2246 2696 2251 2701
rect 2308 2703 2383 2707
rect 2165 2690 2210 2693
rect 2165 2680 2168 2690
rect 2183 2677 2203 2680
rect 2200 2658 2203 2677
rect 2103 2635 2106 2650
rect 2118 2635 2121 2650
rect 2125 2642 2129 2645
rect 2146 2635 2149 2650
rect 1996 2616 1999 2631
rect 2010 2620 2013 2624
rect 2028 2616 2031 2631
rect 2047 2616 2050 2631
rect 1996 2569 1999 2582
rect 2022 2576 2025 2579
rect 1996 2552 1999 2565
rect 2006 2562 2010 2572
rect 2029 2569 2032 2582
rect 2046 2569 2049 2582
rect 2053 2576 2056 2617
rect 2069 2583 2072 2624
rect 2075 2576 2078 2616
rect 2094 2583 2097 2624
rect 2103 2616 2106 2631
rect 2118 2616 2121 2631
rect 2125 2621 2129 2624
rect 2146 2616 2149 2631
rect 2103 2569 2106 2582
rect 2022 2555 2025 2558
rect 2029 2552 2032 2565
rect 2046 2552 2049 2565
rect 1996 2503 1999 2518
rect 2010 2510 2013 2514
rect 2028 2503 2031 2518
rect 2047 2503 2050 2518
rect 2053 2517 2056 2558
rect 2069 2510 2072 2551
rect 2075 2518 2078 2558
rect 2094 2510 2097 2551
rect 2103 2552 2106 2565
rect 2119 2569 2122 2582
rect 2140 2576 2143 2579
rect 2147 2569 2150 2582
rect 2200 2582 2203 2654
rect 2211 2618 2214 2690
rect 2246 2693 2249 2696
rect 2246 2690 2291 2693
rect 2246 2680 2249 2690
rect 2119 2552 2122 2565
rect 2140 2555 2143 2558
rect 2147 2552 2150 2565
rect 2200 2548 2203 2578
rect 2211 2562 2214 2614
rect 2218 2602 2222 2668
rect 2206 2558 2210 2561
rect 2199 2545 2203 2548
rect 2200 2526 2203 2545
rect 2103 2503 2106 2518
rect 2118 2503 2121 2518
rect 2125 2510 2129 2513
rect 2146 2503 2149 2518
rect 1996 2484 1999 2499
rect 2010 2488 2013 2492
rect 2028 2484 2031 2499
rect 2047 2484 2050 2499
rect 1996 2437 1999 2450
rect 2022 2444 2025 2447
rect 1996 2420 1999 2433
rect 2029 2437 2032 2450
rect 2046 2437 2049 2450
rect 2053 2444 2056 2485
rect 2069 2451 2072 2492
rect 2075 2444 2078 2484
rect 2094 2451 2097 2492
rect 2103 2484 2106 2499
rect 2118 2484 2121 2499
rect 2125 2489 2129 2492
rect 2146 2484 2149 2499
rect 2103 2437 2106 2450
rect 2022 2423 2025 2426
rect 2029 2420 2032 2433
rect 2046 2420 2049 2433
rect 1996 2371 1999 2386
rect 2010 2378 2013 2382
rect 2028 2371 2031 2386
rect 2047 2371 2050 2386
rect 2053 2385 2056 2426
rect 2069 2378 2072 2419
rect 2075 2386 2078 2426
rect 2094 2378 2097 2419
rect 2103 2420 2106 2433
rect 2119 2437 2122 2450
rect 2140 2444 2143 2447
rect 2147 2437 2150 2450
rect 2200 2451 2203 2522
rect 2211 2487 2214 2558
rect 2119 2420 2122 2433
rect 2140 2423 2143 2426
rect 2147 2420 2150 2433
rect 2200 2394 2203 2447
rect 2211 2430 2214 2483
rect 2218 2471 2222 2536
rect 2206 2426 2210 2429
rect 2249 2429 2252 2680
rect 2264 2677 2284 2680
rect 2281 2658 2284 2677
rect 2281 2582 2284 2654
rect 2292 2618 2295 2690
rect 2299 2602 2303 2668
rect 2308 2569 2311 2703
rect 2512 2700 2515 2729
rect 2336 2697 2443 2700
rect 2270 2565 2311 2569
rect 2270 2561 2273 2565
rect 2270 2558 2315 2561
rect 2270 2548 2273 2558
rect 2288 2545 2308 2548
rect 2270 2543 2273 2544
rect 2305 2526 2308 2545
rect 2305 2451 2308 2522
rect 2316 2487 2319 2558
rect 2323 2471 2327 2536
rect 2103 2371 2106 2386
rect 2118 2371 2121 2386
rect 2125 2378 2129 2381
rect 2146 2371 2149 2386
rect 1996 2352 1999 2367
rect 2010 2356 2013 2360
rect 2028 2352 2031 2367
rect 2047 2352 2050 2367
rect 1996 2305 1999 2318
rect 2022 2312 2025 2315
rect 1996 2288 1999 2301
rect 2029 2305 2032 2318
rect 2046 2305 2049 2318
rect 2053 2312 2056 2353
rect 2069 2319 2072 2360
rect 2075 2312 2078 2352
rect 2094 2319 2097 2360
rect 2103 2352 2106 2367
rect 2118 2352 2121 2367
rect 2125 2357 2129 2360
rect 2146 2352 2149 2367
rect 2103 2305 2106 2318
rect 2022 2291 2025 2294
rect 2029 2288 2032 2301
rect 2046 2288 2049 2301
rect 1996 2239 1999 2254
rect 2010 2246 2013 2250
rect 1996 2220 1999 2235
rect 2019 2232 2023 2242
rect 2028 2239 2031 2254
rect 2047 2239 2050 2254
rect 2053 2253 2056 2294
rect 2069 2246 2072 2287
rect 2075 2254 2078 2294
rect 2094 2246 2097 2287
rect 2103 2288 2106 2301
rect 2119 2305 2122 2318
rect 2140 2312 2143 2315
rect 2147 2305 2150 2318
rect 2200 2316 2203 2390
rect 2211 2352 2214 2426
rect 2246 2426 2291 2429
rect 2246 2416 2249 2426
rect 2264 2413 2284 2416
rect 2119 2288 2122 2301
rect 2140 2291 2143 2294
rect 2147 2288 2150 2301
rect 2200 2262 2203 2312
rect 2211 2298 2214 2348
rect 2218 2336 2222 2404
rect 2281 2394 2284 2413
rect 2281 2316 2284 2390
rect 2292 2352 2295 2426
rect 2336 2429 2339 2697
rect 2447 2697 2515 2700
rect 2575 2665 2578 2714
rect 2575 2621 2578 2661
rect 2583 2658 2587 3100
rect 2591 3076 2594 3086
rect 2598 3046 2601 3055
rect 2614 3048 2617 3061
rect 2627 3033 2630 3086
rect 2694 3076 2697 3086
rect 2634 3061 2638 3065
rect 2635 3046 2638 3055
rect 2590 3019 2593 3031
rect 2631 3029 2632 3033
rect 2641 3019 2644 3072
rect 2647 3052 2650 3057
rect 2656 3046 2659 3055
rect 2672 3048 2675 3061
rect 2693 3046 2696 3055
rect 2692 3019 2695 3029
rect 2591 2990 2594 3000
rect 2598 2960 2601 2969
rect 2614 2962 2617 2975
rect 2627 2947 2630 3000
rect 2694 2990 2697 3000
rect 2634 2975 2638 2979
rect 2635 2960 2638 2969
rect 2590 2933 2593 2945
rect 2631 2943 2632 2947
rect 2641 2933 2644 2986
rect 2647 2966 2650 2971
rect 2656 2960 2659 2969
rect 2672 2962 2675 2975
rect 2693 2960 2696 2969
rect 2692 2933 2695 2943
rect 2700 2912 2704 3645
rect 2724 3640 2728 3645
rect 2849 3625 2855 3679
rect 2849 3551 2855 3621
rect 2849 3419 2855 3547
rect 2849 3287 2855 3415
rect 2723 3218 2726 3228
rect 2709 3188 2712 3197
rect 2730 3188 2733 3197
rect 2746 3190 2749 3203
rect 2709 3147 2712 3184
rect 2759 3175 2762 3228
rect 2826 3218 2829 3228
rect 2849 3225 2855 3283
rect 2766 3203 2770 3207
rect 2767 3188 2770 3197
rect 2722 3161 2725 3173
rect 2763 3171 2764 3175
rect 2773 3161 2776 3214
rect 2779 3194 2782 3199
rect 2788 3188 2791 3197
rect 2804 3190 2807 3203
rect 2825 3188 2828 3197
rect 2841 3188 2844 3199
rect 2824 3161 2827 3171
rect 2841 3154 2844 3184
rect 2841 3120 2844 3150
rect 2849 3155 2855 3221
rect 2849 3113 2855 3151
rect 2709 3061 2712 3093
rect 2723 3076 2726 3086
rect 2709 3046 2712 3055
rect 2730 3046 2733 3055
rect 2746 3048 2749 3061
rect 2759 3033 2762 3086
rect 2826 3076 2829 3086
rect 2766 3061 2770 3065
rect 2767 3046 2770 3055
rect 2722 3019 2725 3031
rect 2763 3029 2764 3033
rect 2773 3019 2776 3072
rect 2841 3061 2844 3108
rect 2779 3052 2782 3057
rect 2788 3046 2791 3055
rect 2804 3048 2807 3061
rect 2825 3046 2828 3055
rect 2841 3046 2844 3057
rect 2824 3019 2827 3029
rect 2841 3012 2844 3042
rect 2849 3083 2855 3109
rect 2723 2990 2726 3000
rect 2709 2960 2712 2969
rect 2730 2960 2733 2969
rect 2746 2962 2749 2975
rect 2709 2919 2712 2956
rect 2759 2947 2762 3000
rect 2826 2990 2829 3000
rect 2849 2997 2855 3079
rect 2766 2975 2770 2979
rect 2767 2960 2770 2969
rect 2722 2933 2725 2945
rect 2763 2943 2764 2947
rect 2773 2933 2776 2986
rect 2779 2966 2782 2971
rect 2788 2960 2791 2969
rect 2804 2962 2807 2975
rect 2825 2960 2828 2969
rect 2841 2960 2844 2971
rect 2824 2933 2827 2943
rect 2841 2926 2844 2956
rect 2684 2901 2688 2904
rect 2684 2882 2688 2897
rect 2700 2894 2704 2908
rect 2716 2908 2720 2912
rect 2716 2901 2720 2904
rect 2716 2882 2720 2897
rect 2841 2894 2844 2922
rect 2700 2878 2704 2879
rect 2716 2874 2720 2878
rect 2591 2850 2594 2860
rect 2598 2820 2601 2829
rect 2614 2822 2617 2835
rect 2627 2807 2630 2860
rect 2694 2850 2697 2860
rect 2634 2835 2638 2839
rect 2635 2820 2638 2829
rect 2590 2793 2593 2805
rect 2631 2803 2632 2807
rect 2641 2793 2644 2846
rect 2647 2826 2650 2831
rect 2656 2820 2659 2829
rect 2672 2822 2675 2835
rect 2693 2820 2696 2829
rect 2692 2793 2695 2803
rect 2591 2738 2594 2748
rect 2598 2708 2601 2717
rect 2614 2710 2617 2723
rect 2627 2695 2630 2748
rect 2694 2738 2697 2748
rect 2634 2723 2638 2727
rect 2635 2708 2638 2717
rect 2590 2681 2593 2693
rect 2631 2691 2632 2695
rect 2641 2681 2644 2734
rect 2647 2714 2650 2719
rect 2656 2708 2659 2717
rect 2672 2710 2675 2723
rect 2693 2708 2696 2717
rect 2692 2681 2695 2691
rect 2575 2606 2578 2615
rect 2336 2426 2381 2429
rect 2336 2416 2339 2426
rect 2354 2413 2374 2416
rect 2299 2336 2303 2404
rect 2371 2394 2374 2413
rect 2371 2316 2374 2390
rect 2382 2352 2385 2426
rect 2389 2336 2393 2404
rect 2206 2294 2210 2297
rect 2103 2239 2106 2254
rect 2118 2239 2121 2254
rect 2125 2246 2129 2249
rect 2146 2239 2149 2254
rect 2010 2224 2013 2228
rect 2028 2220 2031 2235
rect 2047 2220 2050 2235
rect 1996 2173 1999 2186
rect 2022 2180 2025 2183
rect 2004 2166 2008 2176
rect 2029 2173 2032 2186
rect 2046 2173 2049 2186
rect 2053 2180 2056 2221
rect 2069 2187 2072 2228
rect 2075 2180 2078 2220
rect 2094 2187 2097 2228
rect 2103 2220 2106 2235
rect 2118 2220 2121 2235
rect 2125 2225 2129 2228
rect 2146 2220 2149 2235
rect 2103 2173 2106 2186
rect 2119 2173 2122 2186
rect 2140 2180 2143 2183
rect 2147 2173 2150 2186
rect 2200 2180 2203 2258
rect 2211 2216 2214 2294
rect 2218 2200 2222 2272
rect 2230 2173 2234 2186
rect 2239 2166 2242 2176
rect 2249 2159 2252 2228
rect 2271 2224 2274 2228
rect 2289 2220 2292 2235
rect 2308 2220 2311 2235
rect 2256 2173 2260 2186
rect 2283 2180 2286 2183
rect 2290 2173 2293 2186
rect 2307 2173 2310 2186
rect 2314 2180 2317 2221
rect 2330 2187 2333 2228
rect 2336 2180 2339 2220
rect 2355 2187 2358 2228
rect 2364 2220 2367 2235
rect 2379 2220 2382 2235
rect 2386 2225 2390 2228
rect 2407 2220 2410 2235
rect 2364 2173 2367 2186
rect 2380 2173 2383 2186
rect 2401 2180 2404 2183
rect 2408 2173 2411 2186
rect 2424 2167 2428 2403
rect 2459 2236 2462 2246
rect 2466 2206 2469 2215
rect 2482 2208 2485 2221
rect 2495 2193 2498 2246
rect 2562 2236 2565 2246
rect 2502 2221 2506 2225
rect 2503 2206 2506 2215
rect 2458 2179 2461 2191
rect 2499 2189 2500 2193
rect 2509 2179 2512 2232
rect 2515 2212 2518 2217
rect 2524 2206 2527 2215
rect 2540 2208 2543 2221
rect 2561 2206 2564 2215
rect 2577 2206 2580 2215
rect 2560 2179 2563 2189
rect 2417 2155 2418 2158
rect 1976 1797 1982 2148
rect 2282 2045 2286 2127
rect 2297 2124 2300 2134
rect 2304 2094 2307 2103
rect 2320 2096 2323 2109
rect 2333 2081 2336 2134
rect 2400 2124 2403 2134
rect 2340 2109 2344 2113
rect 2341 2094 2344 2103
rect 2296 2067 2299 2079
rect 2337 2077 2338 2081
rect 2347 2067 2350 2120
rect 2415 2109 2418 2155
rect 2353 2100 2356 2105
rect 2362 2094 2365 2103
rect 2378 2096 2381 2109
rect 2399 2094 2402 2103
rect 2415 2094 2418 2103
rect 2398 2067 2401 2077
rect 2415 2060 2418 2090
rect 2290 2018 2293 2055
rect 2297 2038 2300 2048
rect 2304 2008 2307 2017
rect 2320 2010 2323 2023
rect 2333 1995 2336 2048
rect 2400 2038 2403 2048
rect 2340 2023 2344 2027
rect 2341 2008 2344 2017
rect 2296 1981 2299 1993
rect 2337 1991 2338 1995
rect 2347 1981 2350 2034
rect 2353 2014 2356 2019
rect 2362 2008 2365 2017
rect 2378 2010 2381 2023
rect 2399 2008 2402 2017
rect 2415 2018 2418 2019
rect 2436 2021 2440 2163
rect 2452 2074 2455 2168
rect 2577 2165 2580 2202
rect 2583 2158 2587 2654
rect 2700 2667 2704 2874
rect 2709 2835 2712 2867
rect 2723 2850 2726 2860
rect 2709 2820 2712 2829
rect 2730 2820 2733 2829
rect 2746 2822 2749 2835
rect 2759 2807 2762 2860
rect 2826 2850 2829 2860
rect 2766 2835 2770 2839
rect 2767 2820 2770 2829
rect 2722 2793 2725 2805
rect 2763 2803 2764 2807
rect 2773 2793 2776 2846
rect 2841 2835 2844 2882
rect 2779 2826 2782 2831
rect 2788 2820 2791 2829
rect 2804 2822 2807 2835
rect 2825 2820 2828 2829
rect 2841 2827 2844 2831
rect 2849 2857 2855 2993
rect 2841 2820 2844 2823
rect 2824 2793 2827 2803
rect 2849 2778 2855 2853
rect 2849 2745 2855 2774
rect 2709 2716 2712 2717
rect 2709 2711 2713 2712
rect 2709 2708 2712 2711
rect 2709 2674 2712 2704
rect 2849 2701 2855 2741
rect 2590 2636 2593 2646
rect 2591 2606 2594 2615
rect 2612 2608 2615 2621
rect 2628 2606 2631 2615
rect 2637 2612 2640 2617
rect 2592 2579 2595 2589
rect 2643 2579 2646 2632
rect 2649 2621 2653 2625
rect 2649 2606 2652 2615
rect 2657 2593 2660 2646
rect 2693 2636 2696 2646
rect 2670 2608 2673 2621
rect 2686 2606 2689 2615
rect 2655 2589 2656 2593
rect 2694 2579 2697 2591
rect 2591 2236 2594 2246
rect 2598 2206 2601 2215
rect 2614 2208 2617 2221
rect 2627 2193 2630 2246
rect 2694 2236 2697 2246
rect 2634 2221 2638 2225
rect 2635 2206 2638 2215
rect 2590 2179 2593 2191
rect 2631 2189 2632 2193
rect 2641 2179 2644 2232
rect 2647 2212 2650 2217
rect 2656 2206 2659 2215
rect 2672 2208 2675 2221
rect 2693 2206 2696 2215
rect 2692 2179 2695 2189
rect 2567 2145 2571 2150
rect 2567 2126 2571 2141
rect 2583 2138 2587 2154
rect 2599 2154 2603 2158
rect 2599 2145 2603 2150
rect 2599 2126 2603 2141
rect 2583 2122 2587 2123
rect 2599 2118 2603 2122
rect 2459 2094 2462 2104
rect 2466 2064 2469 2073
rect 2482 2066 2485 2079
rect 2495 2051 2498 2104
rect 2562 2094 2565 2104
rect 2502 2079 2506 2083
rect 2503 2064 2506 2073
rect 2458 2037 2461 2049
rect 2499 2047 2500 2051
rect 2509 2037 2512 2090
rect 2577 2079 2580 2111
rect 2515 2070 2518 2075
rect 2524 2064 2527 2073
rect 2540 2066 2543 2079
rect 2561 2064 2564 2073
rect 2577 2064 2580 2073
rect 2560 2037 2563 2047
rect 2415 2013 2418 2014
rect 2398 1981 2401 1991
rect 2436 1919 2440 2001
rect 2452 1988 2455 2026
rect 2459 2008 2462 2018
rect 2466 1978 2469 1987
rect 2482 1980 2485 1993
rect 2495 1965 2498 2018
rect 2562 2008 2565 2018
rect 2502 1993 2506 1997
rect 2503 1978 2506 1987
rect 2458 1951 2461 1963
rect 2499 1961 2500 1965
rect 2509 1951 2512 2004
rect 2515 1984 2518 1989
rect 2524 1978 2527 1987
rect 2540 1980 2543 1993
rect 2561 1978 2564 1987
rect 2577 1978 2580 1987
rect 2560 1951 2563 1961
rect 2452 1848 2455 1940
rect 2577 1937 2580 1974
rect 2459 1868 2462 1878
rect 2466 1838 2469 1847
rect 2482 1840 2485 1853
rect 2495 1825 2498 1878
rect 2562 1868 2565 1878
rect 2502 1853 2506 1857
rect 2503 1838 2506 1847
rect 2458 1811 2461 1823
rect 2499 1821 2500 1825
rect 2509 1811 2512 1864
rect 2577 1853 2580 1885
rect 2515 1844 2518 1849
rect 2524 1838 2527 1847
rect 2540 1840 2543 1853
rect 2561 1838 2564 1847
rect 2577 1838 2580 1847
rect 2560 1811 2563 1821
rect 2583 1797 2587 2118
rect 2591 2094 2594 2104
rect 2598 2064 2601 2073
rect 2614 2066 2617 2079
rect 2627 2051 2630 2104
rect 2694 2094 2697 2104
rect 2634 2079 2638 2083
rect 2635 2064 2638 2073
rect 2590 2037 2593 2049
rect 2631 2047 2632 2051
rect 2641 2037 2644 2090
rect 2647 2070 2650 2075
rect 2656 2064 2659 2073
rect 2672 2066 2675 2079
rect 2693 2064 2696 2073
rect 2692 2037 2695 2047
rect 2591 2008 2594 2018
rect 2598 1978 2601 1987
rect 2614 1980 2617 1993
rect 2627 1965 2630 2018
rect 2694 2008 2697 2018
rect 2634 1993 2638 1997
rect 2635 1978 2638 1987
rect 2590 1951 2593 1963
rect 2631 1961 2632 1965
rect 2641 1951 2644 2004
rect 2647 1984 2650 1989
rect 2656 1978 2659 1987
rect 2672 1980 2675 1993
rect 2693 1978 2696 1987
rect 2692 1951 2695 1961
rect 2700 1930 2704 2663
rect 2724 2658 2728 2663
rect 2849 2643 2855 2697
rect 2849 2569 2855 2639
rect 2849 2437 2855 2565
rect 2849 2305 2855 2433
rect 2723 2236 2726 2246
rect 2709 2206 2712 2215
rect 2730 2206 2733 2215
rect 2746 2208 2749 2221
rect 2709 2165 2712 2202
rect 2759 2193 2762 2246
rect 2826 2236 2829 2246
rect 2849 2243 2855 2301
rect 2766 2221 2770 2225
rect 2767 2206 2770 2215
rect 2722 2179 2725 2191
rect 2763 2189 2764 2193
rect 2773 2179 2776 2232
rect 2779 2212 2782 2217
rect 2788 2206 2791 2215
rect 2804 2208 2807 2221
rect 2825 2206 2828 2215
rect 2841 2206 2844 2217
rect 2824 2179 2827 2189
rect 2841 2172 2844 2202
rect 2841 2138 2844 2168
rect 2849 2173 2855 2239
rect 2849 2131 2855 2169
rect 2709 2079 2712 2111
rect 2723 2094 2726 2104
rect 2709 2064 2712 2073
rect 2730 2064 2733 2073
rect 2746 2066 2749 2079
rect 2759 2051 2762 2104
rect 2826 2094 2829 2104
rect 2766 2079 2770 2083
rect 2767 2064 2770 2073
rect 2722 2037 2725 2049
rect 2763 2047 2764 2051
rect 2773 2037 2776 2090
rect 2841 2079 2844 2126
rect 2779 2070 2782 2075
rect 2788 2064 2791 2073
rect 2804 2066 2807 2079
rect 2825 2064 2828 2073
rect 2841 2064 2844 2075
rect 2824 2037 2827 2047
rect 2841 2030 2844 2060
rect 2849 2101 2855 2127
rect 2723 2008 2726 2018
rect 2709 1978 2712 1987
rect 2730 1978 2733 1987
rect 2746 1980 2749 1993
rect 2709 1937 2712 1974
rect 2759 1965 2762 2018
rect 2826 2008 2829 2018
rect 2849 2015 2855 2097
rect 2766 1993 2770 1997
rect 2767 1978 2770 1987
rect 2722 1951 2725 1963
rect 2763 1961 2764 1965
rect 2773 1951 2776 2004
rect 2779 1984 2782 1989
rect 2788 1978 2791 1987
rect 2804 1980 2807 1993
rect 2825 1978 2828 1987
rect 2841 1978 2844 1989
rect 2824 1951 2827 1961
rect 2841 1944 2844 1974
rect 2684 1919 2688 1922
rect 2684 1900 2688 1915
rect 2700 1912 2704 1926
rect 2716 1926 2720 1930
rect 2716 1919 2720 1922
rect 2716 1900 2720 1915
rect 2841 1912 2844 1940
rect 2700 1896 2704 1897
rect 2716 1892 2720 1896
rect 2591 1868 2594 1878
rect 2598 1838 2601 1847
rect 2614 1840 2617 1853
rect 2627 1825 2630 1878
rect 2694 1868 2697 1878
rect 2634 1853 2638 1857
rect 2635 1838 2638 1847
rect 2590 1811 2593 1823
rect 2631 1821 2632 1825
rect 2641 1811 2644 1864
rect 2647 1844 2650 1849
rect 2656 1838 2659 1847
rect 2672 1840 2675 1853
rect 2693 1838 2696 1847
rect 2692 1811 2695 1821
rect 2700 1797 2704 1892
rect 2709 1853 2712 1885
rect 2723 1868 2726 1878
rect 2709 1838 2712 1847
rect 2730 1838 2733 1847
rect 2746 1840 2749 1853
rect 2759 1825 2762 1878
rect 2826 1868 2829 1878
rect 2766 1853 2770 1857
rect 2767 1838 2770 1847
rect 2722 1811 2725 1823
rect 2763 1821 2764 1825
rect 2773 1811 2776 1864
rect 2841 1853 2844 1900
rect 2779 1844 2782 1849
rect 2788 1838 2791 1847
rect 2804 1840 2807 1853
rect 2825 1838 2828 1847
rect 2841 1845 2844 1849
rect 2849 1875 2855 2011
rect 2841 1838 2844 1841
rect 2824 1811 2827 1821
rect 2849 1797 2855 1871
rect 2861 3816 2867 3921
rect 2861 3808 2867 3812
rect 2861 3703 2867 3804
rect 2861 3670 2867 3699
rect 2861 3617 2867 3666
rect 2861 3568 2867 3613
rect 2861 3485 2867 3564
rect 2861 3353 2867 3481
rect 2861 3221 2867 3349
rect 2861 3168 2867 3217
rect 2861 3056 2867 3164
rect 2861 3026 2867 3052
rect 2861 2970 2867 3022
rect 2861 2940 2867 2966
rect 2861 2800 2867 2936
rect 2861 2721 2867 2796
rect 2861 2688 2867 2717
rect 2861 2635 2867 2684
rect 2861 2586 2867 2631
rect 2861 2503 2867 2582
rect 2861 2371 2867 2499
rect 2861 2239 2867 2367
rect 2861 2186 2867 2235
rect 2861 2074 2867 2182
rect 2861 2044 2867 2070
rect 2861 1988 2867 2040
rect 2861 1958 2867 1984
rect 2861 1818 2867 1954
rect 2861 1797 2867 1814
rect 2873 3932 2879 3987
rect 2873 3824 2879 3928
rect 2873 3816 2879 3820
rect 2873 3624 2879 3812
rect 2873 3610 2879 3620
rect 2873 3492 2879 3606
rect 2873 3478 2879 3488
rect 2873 3360 2879 3474
rect 2873 3346 2879 3356
rect 2873 3214 2879 3342
rect 2873 3140 2879 3210
rect 2873 2642 2879 3136
rect 2873 2628 2879 2638
rect 2873 2510 2879 2624
rect 2873 2496 2879 2506
rect 2873 2378 2879 2492
rect 2873 2364 2879 2374
rect 2873 2232 2879 2360
rect 2873 2158 2879 2228
rect 2873 1797 2879 2154
rect 2885 3939 2891 4059
rect 2885 3832 2891 3935
rect 2885 3824 2891 3828
rect 2885 3676 2891 3820
rect 2885 3544 2891 3672
rect 2885 3426 2891 3540
rect 2885 3412 2891 3422
rect 2885 3294 2891 3408
rect 2885 3280 2891 3290
rect 2885 3148 2891 3276
rect 2885 2694 2891 3144
rect 2885 2562 2891 2690
rect 2885 2444 2891 2558
rect 2885 2430 2891 2440
rect 2885 2312 2891 2426
rect 2885 2298 2891 2308
rect 2885 2166 2891 2294
rect 2885 1797 2891 2162
rect 2897 3947 2903 4102
rect 2923 3998 2927 4231
rect 2956 4204 2960 4231
rect 2930 4200 2960 4204
rect 2990 4204 2995 4294
rect 2930 3991 2934 4200
rect 2990 4074 2995 4200
rect 2897 3840 2903 3943
rect 2990 3917 2995 4070
rect 2998 4154 3002 4264
rect 2998 4024 3002 4150
rect 2998 3910 3002 4020
rect 3006 3902 3010 4246
rect 2897 3832 2903 3836
rect 2897 3696 2903 3828
rect 2897 3663 2903 3692
rect 2897 3561 2903 3659
rect 2897 3162 2903 3557
rect 2897 3049 2903 3158
rect 2897 3019 2903 3045
rect 2897 2963 2903 3015
rect 2897 2933 2903 2959
rect 2897 2793 2903 2929
rect 2897 2714 2903 2789
rect 2897 2681 2903 2710
rect 2897 2579 2903 2677
rect 2897 2180 2903 2575
rect 2897 2067 2903 2176
rect 2897 2037 2903 2063
rect 2897 1981 2903 2033
rect 2897 1951 2903 1977
rect 2897 1811 2903 1947
rect 2897 1797 2903 1807
rect 2909 3767 2915 3836
rect 2909 3734 2915 3763
rect 2909 3632 2915 3730
rect 2909 3232 2915 3628
rect 2909 3120 2915 3228
rect 2909 3090 2915 3116
rect 2909 3034 2915 3086
rect 2909 3004 2915 3030
rect 2909 2864 2915 3000
rect 2909 2785 2915 2860
rect 2909 2752 2915 2781
rect 2909 2650 2915 2748
rect 2909 2250 2915 2646
rect 2909 2138 2915 2246
rect 2909 2108 2915 2134
rect 2909 2052 2915 2104
rect 2909 2022 2915 2048
rect 2909 1882 2915 2018
rect 2909 1797 2915 1878
rect 2921 3134 2927 3898
rect 2943 3753 2946 3763
rect 2950 3723 2953 3732
rect 2966 3725 2969 3738
rect 2979 3710 2982 3763
rect 3046 3753 3049 3763
rect 3075 3753 3078 3763
rect 2986 3738 2990 3742
rect 2987 3723 2990 3732
rect 2942 3696 2945 3708
rect 2983 3706 2984 3710
rect 2993 3696 2996 3749
rect 2999 3729 3002 3734
rect 3008 3723 3011 3732
rect 3024 3725 3027 3738
rect 3045 3723 3048 3732
rect 3061 3732 3064 3734
rect 3061 3729 3068 3732
rect 3061 3723 3064 3729
rect 3082 3723 3085 3732
rect 3098 3725 3101 3738
rect 3044 3696 3047 3706
rect 3061 3689 3064 3719
rect 3111 3710 3114 3763
rect 3178 3753 3181 3763
rect 3207 3753 3210 3763
rect 3118 3738 3122 3742
rect 3119 3723 3122 3732
rect 3074 3696 3077 3708
rect 3115 3706 3116 3710
rect 3125 3696 3128 3749
rect 3131 3729 3134 3734
rect 3140 3723 3143 3732
rect 3156 3725 3159 3738
rect 3177 3723 3180 3732
rect 3193 3732 3196 3734
rect 3193 3729 3200 3732
rect 3193 3723 3196 3729
rect 3214 3723 3217 3732
rect 3230 3725 3233 3738
rect 3176 3696 3179 3706
rect 3061 3686 3113 3689
rect 2941 3666 2944 3679
rect 2967 3669 2970 3672
rect 2974 3666 2977 3679
rect 2991 3666 2994 3679
rect 2941 3617 2944 3632
rect 2955 3624 2958 3628
rect 2973 3617 2976 3632
rect 2992 3617 2995 3632
rect 2998 3631 3001 3672
rect 3014 3624 3017 3665
rect 3020 3632 3023 3672
rect 3039 3624 3042 3665
rect 3048 3666 3051 3679
rect 3064 3666 3067 3679
rect 3085 3669 3088 3672
rect 3092 3666 3095 3679
rect 3110 3675 3113 3686
rect 3193 3683 3196 3719
rect 3243 3710 3246 3763
rect 3310 3753 3313 3763
rect 3339 3753 3342 3763
rect 3250 3738 3254 3742
rect 3251 3723 3254 3732
rect 3206 3696 3209 3708
rect 3247 3706 3248 3710
rect 3257 3696 3260 3749
rect 3263 3729 3266 3734
rect 3272 3723 3275 3732
rect 3288 3725 3291 3738
rect 3309 3723 3312 3732
rect 3325 3732 3328 3734
rect 3325 3729 3332 3732
rect 3325 3723 3328 3729
rect 3346 3723 3349 3732
rect 3362 3725 3365 3738
rect 3308 3696 3311 3706
rect 3325 3689 3328 3711
rect 3375 3710 3378 3763
rect 3442 3753 3445 3763
rect 3382 3738 3386 3742
rect 3383 3723 3386 3732
rect 3338 3696 3341 3708
rect 3379 3706 3380 3710
rect 3389 3696 3392 3749
rect 3395 3729 3398 3734
rect 3404 3723 3407 3732
rect 3420 3725 3423 3738
rect 3441 3723 3444 3732
rect 3457 3732 3460 3734
rect 3457 3729 3461 3732
rect 3457 3723 3460 3729
rect 3457 3715 3460 3719
rect 3440 3696 3443 3706
rect 3191 3678 3196 3683
rect 3253 3685 3328 3689
rect 3110 3672 3155 3675
rect 3110 3662 3113 3672
rect 3128 3659 3148 3662
rect 3145 3640 3148 3659
rect 3048 3617 3051 3632
rect 3063 3617 3066 3632
rect 3070 3624 3074 3627
rect 3091 3617 3094 3632
rect 2941 3598 2944 3613
rect 2955 3602 2958 3606
rect 2973 3598 2976 3613
rect 2992 3598 2995 3613
rect 2941 3551 2944 3564
rect 2967 3558 2970 3561
rect 2941 3534 2944 3547
rect 2951 3544 2955 3554
rect 2974 3551 2977 3564
rect 2991 3551 2994 3564
rect 2998 3558 3001 3599
rect 3014 3565 3017 3606
rect 3020 3558 3023 3598
rect 3039 3565 3042 3606
rect 3048 3598 3051 3613
rect 3063 3598 3066 3613
rect 3070 3603 3074 3606
rect 3091 3598 3094 3613
rect 3048 3551 3051 3564
rect 2967 3537 2970 3540
rect 2974 3534 2977 3547
rect 2991 3534 2994 3547
rect 2941 3485 2944 3500
rect 2955 3492 2958 3496
rect 2973 3485 2976 3500
rect 2992 3485 2995 3500
rect 2998 3499 3001 3540
rect 3014 3492 3017 3533
rect 3020 3500 3023 3540
rect 3039 3492 3042 3533
rect 3048 3534 3051 3547
rect 3064 3551 3067 3564
rect 3085 3558 3088 3561
rect 3092 3551 3095 3564
rect 3145 3564 3148 3636
rect 3156 3600 3159 3672
rect 3191 3675 3194 3678
rect 3191 3672 3236 3675
rect 3191 3662 3194 3672
rect 3064 3534 3067 3547
rect 3085 3537 3088 3540
rect 3092 3534 3095 3547
rect 3145 3530 3148 3560
rect 3156 3544 3159 3596
rect 3163 3584 3167 3650
rect 3151 3540 3155 3543
rect 3144 3527 3148 3530
rect 3145 3508 3148 3527
rect 3048 3485 3051 3500
rect 3063 3485 3066 3500
rect 3070 3492 3074 3495
rect 3091 3485 3094 3500
rect 2941 3466 2944 3481
rect 2955 3470 2958 3474
rect 2973 3466 2976 3481
rect 2992 3466 2995 3481
rect 2941 3419 2944 3432
rect 2967 3426 2970 3429
rect 2941 3402 2944 3415
rect 2974 3419 2977 3432
rect 2991 3419 2994 3432
rect 2998 3426 3001 3467
rect 3014 3433 3017 3474
rect 3020 3426 3023 3466
rect 3039 3433 3042 3474
rect 3048 3466 3051 3481
rect 3063 3466 3066 3481
rect 3070 3471 3074 3474
rect 3091 3466 3094 3481
rect 3048 3419 3051 3432
rect 2967 3405 2970 3408
rect 2974 3402 2977 3415
rect 2991 3402 2994 3415
rect 2941 3353 2944 3368
rect 2955 3360 2958 3364
rect 2973 3353 2976 3368
rect 2992 3353 2995 3368
rect 2998 3367 3001 3408
rect 3014 3360 3017 3401
rect 3020 3368 3023 3408
rect 3039 3360 3042 3401
rect 3048 3402 3051 3415
rect 3064 3419 3067 3432
rect 3085 3426 3088 3429
rect 3092 3419 3095 3432
rect 3145 3433 3148 3504
rect 3156 3469 3159 3540
rect 3064 3402 3067 3415
rect 3085 3405 3088 3408
rect 3092 3402 3095 3415
rect 3145 3376 3148 3429
rect 3156 3412 3159 3465
rect 3163 3453 3167 3518
rect 3151 3408 3155 3411
rect 3194 3411 3197 3662
rect 3209 3659 3229 3662
rect 3226 3640 3229 3659
rect 3226 3564 3229 3636
rect 3237 3600 3240 3672
rect 3244 3584 3248 3650
rect 3253 3551 3256 3685
rect 3457 3682 3460 3711
rect 3281 3679 3388 3682
rect 3215 3547 3256 3551
rect 3215 3543 3218 3547
rect 3215 3540 3260 3543
rect 3215 3530 3218 3540
rect 3233 3527 3253 3530
rect 3215 3525 3218 3526
rect 3250 3508 3253 3527
rect 3250 3433 3253 3504
rect 3261 3469 3264 3540
rect 3268 3453 3272 3518
rect 3048 3353 3051 3368
rect 3063 3353 3066 3368
rect 3070 3360 3074 3363
rect 3091 3353 3094 3368
rect 2941 3334 2944 3349
rect 2955 3338 2958 3342
rect 2973 3334 2976 3349
rect 2992 3334 2995 3349
rect 2941 3287 2944 3300
rect 2967 3294 2970 3297
rect 2941 3270 2944 3283
rect 2974 3287 2977 3300
rect 2991 3287 2994 3300
rect 2998 3294 3001 3335
rect 3014 3301 3017 3342
rect 3020 3294 3023 3334
rect 3039 3301 3042 3342
rect 3048 3334 3051 3349
rect 3063 3334 3066 3349
rect 3070 3339 3074 3342
rect 3091 3334 3094 3349
rect 3048 3287 3051 3300
rect 2967 3273 2970 3276
rect 2974 3270 2977 3283
rect 2991 3270 2994 3283
rect 2941 3221 2944 3236
rect 2955 3228 2958 3232
rect 2941 3202 2944 3217
rect 2964 3214 2968 3224
rect 2973 3221 2976 3236
rect 2992 3221 2995 3236
rect 2998 3235 3001 3276
rect 3014 3228 3017 3269
rect 3020 3236 3023 3276
rect 3039 3228 3042 3269
rect 3048 3270 3051 3283
rect 3064 3287 3067 3300
rect 3085 3294 3088 3297
rect 3092 3287 3095 3300
rect 3145 3298 3148 3372
rect 3156 3334 3159 3408
rect 3191 3408 3236 3411
rect 3191 3398 3194 3408
rect 3209 3395 3229 3398
rect 3064 3270 3067 3283
rect 3085 3273 3088 3276
rect 3092 3270 3095 3283
rect 3145 3244 3148 3294
rect 3156 3280 3159 3330
rect 3163 3318 3167 3386
rect 3226 3376 3229 3395
rect 3226 3298 3229 3372
rect 3237 3334 3240 3408
rect 3281 3411 3284 3679
rect 3392 3679 3460 3682
rect 3281 3408 3326 3411
rect 3281 3398 3284 3408
rect 3299 3395 3319 3398
rect 3244 3318 3248 3386
rect 3316 3376 3319 3395
rect 3316 3298 3319 3372
rect 3327 3334 3330 3408
rect 3334 3318 3338 3386
rect 3151 3276 3155 3279
rect 3048 3221 3051 3236
rect 3063 3221 3066 3236
rect 3070 3228 3074 3231
rect 3091 3221 3094 3236
rect 2955 3206 2958 3210
rect 2973 3202 2976 3217
rect 2992 3202 2995 3217
rect 2941 3155 2944 3168
rect 2967 3162 2970 3165
rect 2949 3148 2953 3158
rect 2974 3155 2977 3168
rect 2991 3155 2994 3168
rect 2998 3162 3001 3203
rect 3014 3169 3017 3210
rect 3020 3162 3023 3202
rect 3039 3169 3042 3210
rect 3048 3202 3051 3217
rect 3063 3202 3066 3217
rect 3070 3207 3074 3210
rect 3091 3202 3094 3217
rect 3048 3155 3051 3168
rect 3064 3155 3067 3168
rect 3085 3162 3088 3165
rect 3092 3155 3095 3168
rect 3145 3162 3148 3240
rect 3156 3198 3159 3276
rect 3163 3182 3167 3254
rect 3175 3155 3179 3168
rect 3184 3148 3187 3158
rect 3194 3141 3197 3210
rect 3216 3206 3219 3210
rect 3234 3202 3237 3217
rect 3253 3202 3256 3217
rect 3201 3155 3205 3168
rect 3228 3162 3231 3165
rect 3235 3155 3238 3168
rect 3252 3155 3255 3168
rect 3259 3162 3262 3203
rect 3275 3169 3278 3210
rect 3281 3162 3284 3202
rect 3300 3169 3303 3210
rect 3309 3202 3312 3217
rect 3324 3202 3327 3217
rect 3331 3207 3335 3210
rect 3352 3202 3355 3217
rect 3309 3155 3312 3168
rect 3325 3155 3328 3168
rect 3346 3162 3349 3165
rect 3353 3155 3356 3168
rect 3369 3149 3373 3385
rect 3362 3137 3363 3140
rect 2921 2152 2927 3130
rect 3227 3027 3231 3109
rect 3242 3106 3245 3116
rect 3249 3076 3252 3085
rect 3265 3078 3268 3091
rect 3278 3063 3281 3116
rect 3345 3106 3348 3116
rect 3285 3091 3289 3095
rect 3286 3076 3289 3085
rect 3241 3049 3244 3061
rect 3282 3059 3283 3063
rect 3292 3049 3295 3102
rect 3360 3091 3363 3137
rect 3298 3082 3301 3087
rect 3307 3076 3310 3085
rect 3323 3078 3326 3091
rect 3344 3076 3347 3085
rect 3360 3076 3363 3085
rect 3343 3049 3346 3059
rect 3360 3042 3363 3072
rect 3235 3000 3238 3037
rect 3242 3020 3245 3030
rect 3249 2990 3252 2999
rect 3265 2992 3268 3005
rect 3278 2977 3281 3030
rect 3345 3020 3348 3030
rect 3285 3005 3289 3009
rect 3286 2990 3289 2999
rect 3241 2963 3244 2975
rect 3282 2973 3283 2977
rect 3292 2963 3295 3016
rect 3298 2996 3301 3001
rect 3307 2990 3310 2999
rect 3323 2992 3326 3005
rect 3344 2990 3347 2999
rect 3360 3000 3363 3001
rect 3381 3003 3385 3145
rect 3360 2995 3363 2996
rect 3343 2963 3346 2973
rect 3381 2901 3385 2983
rect 2943 2771 2946 2781
rect 2950 2741 2953 2750
rect 2966 2743 2969 2756
rect 2979 2728 2982 2781
rect 3046 2771 3049 2781
rect 3075 2771 3078 2781
rect 2986 2756 2990 2760
rect 2987 2741 2990 2750
rect 2942 2714 2945 2726
rect 2983 2724 2984 2728
rect 2993 2714 2996 2767
rect 2999 2747 3002 2752
rect 3008 2741 3011 2750
rect 3024 2743 3027 2756
rect 3045 2741 3048 2750
rect 3061 2750 3064 2752
rect 3061 2747 3068 2750
rect 3061 2741 3064 2747
rect 3082 2741 3085 2750
rect 3098 2743 3101 2756
rect 3044 2714 3047 2724
rect 3061 2707 3064 2737
rect 3111 2728 3114 2781
rect 3178 2771 3181 2781
rect 3207 2771 3210 2781
rect 3118 2756 3122 2760
rect 3119 2741 3122 2750
rect 3074 2714 3077 2726
rect 3115 2724 3116 2728
rect 3125 2714 3128 2767
rect 3131 2747 3134 2752
rect 3140 2741 3143 2750
rect 3156 2743 3159 2756
rect 3177 2741 3180 2750
rect 3193 2750 3196 2752
rect 3193 2747 3200 2750
rect 3193 2741 3196 2747
rect 3214 2741 3217 2750
rect 3230 2743 3233 2756
rect 3176 2714 3179 2724
rect 3061 2704 3113 2707
rect 2941 2684 2944 2697
rect 2967 2687 2970 2690
rect 2974 2684 2977 2697
rect 2991 2684 2994 2697
rect 2941 2635 2944 2650
rect 2955 2642 2958 2646
rect 2973 2635 2976 2650
rect 2992 2635 2995 2650
rect 2998 2649 3001 2690
rect 3014 2642 3017 2683
rect 3020 2650 3023 2690
rect 3039 2642 3042 2683
rect 3048 2684 3051 2697
rect 3064 2684 3067 2697
rect 3085 2687 3088 2690
rect 3092 2684 3095 2697
rect 3110 2693 3113 2704
rect 3193 2701 3196 2737
rect 3243 2728 3246 2781
rect 3310 2771 3313 2781
rect 3339 2771 3342 2781
rect 3250 2756 3254 2760
rect 3251 2741 3254 2750
rect 3206 2714 3209 2726
rect 3247 2724 3248 2728
rect 3257 2714 3260 2767
rect 3263 2747 3266 2752
rect 3272 2741 3275 2750
rect 3288 2743 3291 2756
rect 3309 2741 3312 2750
rect 3325 2750 3328 2752
rect 3325 2747 3332 2750
rect 3325 2741 3328 2747
rect 3346 2741 3349 2750
rect 3362 2743 3365 2756
rect 3308 2714 3311 2724
rect 3325 2707 3328 2729
rect 3375 2728 3378 2781
rect 3442 2771 3445 2781
rect 3382 2756 3386 2760
rect 3383 2741 3386 2750
rect 3338 2714 3341 2726
rect 3379 2724 3380 2728
rect 3389 2714 3392 2767
rect 3395 2747 3398 2752
rect 3404 2741 3407 2750
rect 3420 2743 3423 2756
rect 3441 2741 3444 2750
rect 3457 2750 3460 2752
rect 3457 2747 3461 2750
rect 3457 2741 3460 2747
rect 3457 2733 3460 2737
rect 3440 2714 3443 2724
rect 3191 2696 3196 2701
rect 3253 2703 3328 2707
rect 3110 2690 3155 2693
rect 3110 2680 3113 2690
rect 3128 2677 3148 2680
rect 3145 2658 3148 2677
rect 3048 2635 3051 2650
rect 3063 2635 3066 2650
rect 3070 2642 3074 2645
rect 3091 2635 3094 2650
rect 2941 2616 2944 2631
rect 2955 2620 2958 2624
rect 2973 2616 2976 2631
rect 2992 2616 2995 2631
rect 2941 2569 2944 2582
rect 2967 2576 2970 2579
rect 2941 2552 2944 2565
rect 2951 2562 2955 2572
rect 2974 2569 2977 2582
rect 2991 2569 2994 2582
rect 2998 2576 3001 2617
rect 3014 2583 3017 2624
rect 3020 2576 3023 2616
rect 3039 2583 3042 2624
rect 3048 2616 3051 2631
rect 3063 2616 3066 2631
rect 3070 2621 3074 2624
rect 3091 2616 3094 2631
rect 3048 2569 3051 2582
rect 2967 2555 2970 2558
rect 2974 2552 2977 2565
rect 2991 2552 2994 2565
rect 2941 2503 2944 2518
rect 2955 2510 2958 2514
rect 2973 2503 2976 2518
rect 2992 2503 2995 2518
rect 2998 2517 3001 2558
rect 3014 2510 3017 2551
rect 3020 2518 3023 2558
rect 3039 2510 3042 2551
rect 3048 2552 3051 2565
rect 3064 2569 3067 2582
rect 3085 2576 3088 2579
rect 3092 2569 3095 2582
rect 3145 2582 3148 2654
rect 3156 2618 3159 2690
rect 3191 2693 3194 2696
rect 3191 2690 3236 2693
rect 3191 2680 3194 2690
rect 3064 2552 3067 2565
rect 3085 2555 3088 2558
rect 3092 2552 3095 2565
rect 3145 2548 3148 2578
rect 3156 2562 3159 2614
rect 3163 2602 3167 2668
rect 3151 2558 3155 2561
rect 3144 2545 3148 2548
rect 3145 2526 3148 2545
rect 3048 2503 3051 2518
rect 3063 2503 3066 2518
rect 3070 2510 3074 2513
rect 3091 2503 3094 2518
rect 2941 2484 2944 2499
rect 2955 2488 2958 2492
rect 2973 2484 2976 2499
rect 2992 2484 2995 2499
rect 2941 2437 2944 2450
rect 2967 2444 2970 2447
rect 2941 2420 2944 2433
rect 2974 2437 2977 2450
rect 2991 2437 2994 2450
rect 2998 2444 3001 2485
rect 3014 2451 3017 2492
rect 3020 2444 3023 2484
rect 3039 2451 3042 2492
rect 3048 2484 3051 2499
rect 3063 2484 3066 2499
rect 3070 2489 3074 2492
rect 3091 2484 3094 2499
rect 3048 2437 3051 2450
rect 2967 2423 2970 2426
rect 2974 2420 2977 2433
rect 2991 2420 2994 2433
rect 2941 2371 2944 2386
rect 2955 2378 2958 2382
rect 2973 2371 2976 2386
rect 2992 2371 2995 2386
rect 2998 2385 3001 2426
rect 3014 2378 3017 2419
rect 3020 2386 3023 2426
rect 3039 2378 3042 2419
rect 3048 2420 3051 2433
rect 3064 2437 3067 2450
rect 3085 2444 3088 2447
rect 3092 2437 3095 2450
rect 3145 2451 3148 2522
rect 3156 2487 3159 2558
rect 3064 2420 3067 2433
rect 3085 2423 3088 2426
rect 3092 2420 3095 2433
rect 3145 2394 3148 2447
rect 3156 2430 3159 2483
rect 3163 2471 3167 2536
rect 3151 2426 3155 2429
rect 3194 2429 3197 2680
rect 3209 2677 3229 2680
rect 3226 2658 3229 2677
rect 3226 2582 3229 2654
rect 3237 2618 3240 2690
rect 3244 2602 3248 2668
rect 3253 2569 3256 2703
rect 3457 2700 3460 2729
rect 3281 2697 3388 2700
rect 3215 2565 3256 2569
rect 3215 2561 3218 2565
rect 3215 2558 3260 2561
rect 3215 2548 3218 2558
rect 3233 2545 3253 2548
rect 3215 2543 3218 2544
rect 3250 2526 3253 2545
rect 3250 2451 3253 2522
rect 3261 2487 3264 2558
rect 3268 2471 3272 2536
rect 3048 2371 3051 2386
rect 3063 2371 3066 2386
rect 3070 2378 3074 2381
rect 3091 2371 3094 2386
rect 2941 2352 2944 2367
rect 2955 2356 2958 2360
rect 2973 2352 2976 2367
rect 2992 2352 2995 2367
rect 2941 2305 2944 2318
rect 2967 2312 2970 2315
rect 2941 2288 2944 2301
rect 2974 2305 2977 2318
rect 2991 2305 2994 2318
rect 2998 2312 3001 2353
rect 3014 2319 3017 2360
rect 3020 2312 3023 2352
rect 3039 2319 3042 2360
rect 3048 2352 3051 2367
rect 3063 2352 3066 2367
rect 3070 2357 3074 2360
rect 3091 2352 3094 2367
rect 3048 2305 3051 2318
rect 2967 2291 2970 2294
rect 2974 2288 2977 2301
rect 2991 2288 2994 2301
rect 2941 2239 2944 2254
rect 2955 2246 2958 2250
rect 2941 2220 2944 2235
rect 2964 2232 2968 2242
rect 2973 2239 2976 2254
rect 2992 2239 2995 2254
rect 2998 2253 3001 2294
rect 3014 2246 3017 2287
rect 3020 2254 3023 2294
rect 3039 2246 3042 2287
rect 3048 2288 3051 2301
rect 3064 2305 3067 2318
rect 3085 2312 3088 2315
rect 3092 2305 3095 2318
rect 3145 2316 3148 2390
rect 3156 2352 3159 2426
rect 3191 2426 3236 2429
rect 3191 2416 3194 2426
rect 3209 2413 3229 2416
rect 3064 2288 3067 2301
rect 3085 2291 3088 2294
rect 3092 2288 3095 2301
rect 3145 2262 3148 2312
rect 3156 2298 3159 2348
rect 3163 2336 3167 2404
rect 3226 2394 3229 2413
rect 3226 2316 3229 2390
rect 3237 2352 3240 2426
rect 3281 2429 3284 2697
rect 3392 2697 3460 2700
rect 3281 2426 3326 2429
rect 3281 2416 3284 2426
rect 3299 2413 3319 2416
rect 3244 2336 3248 2404
rect 3316 2394 3319 2413
rect 3316 2316 3319 2390
rect 3327 2352 3330 2426
rect 3334 2336 3338 2404
rect 3151 2294 3155 2297
rect 3048 2239 3051 2254
rect 3063 2239 3066 2254
rect 3070 2246 3074 2249
rect 3091 2239 3094 2254
rect 2955 2224 2958 2228
rect 2973 2220 2976 2235
rect 2992 2220 2995 2235
rect 2941 2173 2944 2186
rect 2967 2180 2970 2183
rect 2949 2166 2953 2176
rect 2974 2173 2977 2186
rect 2991 2173 2994 2186
rect 2998 2180 3001 2221
rect 3014 2187 3017 2228
rect 3020 2180 3023 2220
rect 3039 2187 3042 2228
rect 3048 2220 3051 2235
rect 3063 2220 3066 2235
rect 3070 2225 3074 2228
rect 3091 2220 3094 2235
rect 3048 2173 3051 2186
rect 3064 2173 3067 2186
rect 3085 2180 3088 2183
rect 3092 2173 3095 2186
rect 3145 2180 3148 2258
rect 3156 2216 3159 2294
rect 3163 2200 3167 2272
rect 3175 2173 3179 2186
rect 3184 2166 3187 2176
rect 3194 2159 3197 2228
rect 3216 2224 3219 2228
rect 3234 2220 3237 2235
rect 3253 2220 3256 2235
rect 3201 2173 3205 2186
rect 3228 2180 3231 2183
rect 3235 2173 3238 2186
rect 3252 2173 3255 2186
rect 3259 2180 3262 2221
rect 3275 2187 3278 2228
rect 3281 2180 3284 2220
rect 3300 2187 3303 2228
rect 3309 2220 3312 2235
rect 3324 2220 3327 2235
rect 3331 2225 3335 2228
rect 3352 2220 3355 2235
rect 3309 2173 3312 2186
rect 3325 2173 3328 2186
rect 3346 2180 3349 2183
rect 3353 2173 3356 2186
rect 3369 2167 3373 2403
rect 4228 2355 4240 2403
rect 3362 2155 3363 2158
rect 2921 1797 2927 2148
rect 3227 2045 3231 2127
rect 3242 2124 3245 2134
rect 3249 2094 3252 2103
rect 3265 2096 3268 2109
rect 3278 2081 3281 2134
rect 3345 2124 3348 2134
rect 3285 2109 3289 2113
rect 3286 2094 3289 2103
rect 3241 2067 3244 2079
rect 3282 2077 3283 2081
rect 3292 2067 3295 2120
rect 3360 2109 3363 2155
rect 3298 2100 3301 2105
rect 3307 2094 3310 2103
rect 3323 2096 3326 2109
rect 3344 2094 3347 2103
rect 3360 2094 3363 2103
rect 3343 2067 3346 2077
rect 3360 2060 3363 2090
rect 3235 2018 3238 2055
rect 3242 2038 3245 2048
rect 3249 2008 3252 2017
rect 3265 2010 3268 2023
rect 3278 1995 3281 2048
rect 3345 2038 3348 2048
rect 3285 2023 3289 2027
rect 3286 2008 3289 2017
rect 3241 1981 3244 1993
rect 3282 1991 3283 1995
rect 3292 1981 3295 2034
rect 3298 2014 3301 2019
rect 3307 2008 3310 2017
rect 3323 2010 3326 2023
rect 3344 2008 3347 2017
rect 3360 2018 3363 2019
rect 3381 2021 3385 2163
rect 3360 2013 3363 2014
rect 3343 1981 3346 1991
rect 3381 1919 3385 2001
<< m3contact >>
rect 2081 4443 2086 4448
rect 2172 4326 2176 4330
rect 1507 3190 1511 3194
rect 1764 3693 1768 3697
rect 1763 3590 1767 3594
rect 1507 2208 1511 2212
rect 1896 2823 1900 2827
rect 1764 2711 1768 2715
rect 1763 2608 1767 2612
rect 1896 1841 1900 1845
rect 1987 3729 1991 3733
rect 2027 3646 2032 3651
rect 2038 3642 2043 3647
rect 2061 3651 2066 3656
rect 2085 3646 2090 3651
rect 2100 3650 2105 3656
rect 2130 3646 2135 3651
rect 2159 3645 2164 3650
rect 2114 3640 2119 3645
rect 2143 3640 2147 3645
rect 2185 3639 2190 3644
rect 1991 3586 1996 3591
rect 2027 3579 2032 3584
rect 2038 3583 2043 3588
rect 2061 3574 2066 3579
rect 2085 3579 2090 3584
rect 2114 3585 2119 3590
rect 2143 3585 2147 3590
rect 2100 3574 2105 3580
rect 2130 3579 2135 3584
rect 2159 3580 2164 3585
rect 2185 3580 2190 3585
rect 1990 3517 1995 3522
rect 2027 3514 2032 3519
rect 2038 3510 2043 3515
rect 2061 3519 2066 3524
rect 2085 3514 2090 3519
rect 2241 3645 2246 3650
rect 2100 3518 2105 3524
rect 2130 3514 2135 3519
rect 2159 3513 2164 3518
rect 2114 3508 2119 3513
rect 2143 3508 2147 3513
rect 2185 3507 2190 3512
rect 1991 3454 1996 3459
rect 2027 3447 2032 3452
rect 2038 3451 2043 3456
rect 2061 3442 2066 3447
rect 2085 3447 2090 3452
rect 2114 3453 2119 3458
rect 2143 3453 2147 3458
rect 2100 3442 2105 3448
rect 2130 3447 2135 3452
rect 2159 3448 2164 3453
rect 2184 3449 2189 3454
rect 1990 3385 1995 3390
rect 2027 3382 2032 3387
rect 2038 3378 2043 3383
rect 2061 3387 2066 3392
rect 2085 3382 2090 3387
rect 2100 3386 2105 3392
rect 2130 3382 2135 3387
rect 2159 3381 2164 3386
rect 2114 3376 2119 3381
rect 2143 3376 2147 3381
rect 2185 3375 2190 3380
rect 2241 3521 2246 3526
rect 2266 3639 2271 3644
rect 2265 3580 2270 3585
rect 2326 3645 2331 3650
rect 2290 3507 2295 3512
rect 2290 3449 2295 3454
rect 1991 3322 1996 3327
rect 2027 3315 2032 3320
rect 2038 3319 2043 3324
rect 2061 3310 2066 3315
rect 2085 3315 2090 3320
rect 2114 3321 2119 3326
rect 2143 3321 2147 3326
rect 2100 3310 2105 3316
rect 2130 3315 2135 3320
rect 2159 3316 2164 3321
rect 2185 3314 2190 3319
rect 1990 3253 1995 3258
rect 2027 3250 2032 3255
rect 2038 3246 2043 3251
rect 2061 3255 2066 3260
rect 2085 3250 2090 3255
rect 2100 3254 2105 3260
rect 2130 3250 2135 3255
rect 2159 3249 2164 3254
rect 2114 3244 2119 3249
rect 2143 3244 2147 3249
rect 2185 3243 2190 3248
rect 2241 3381 2246 3386
rect 2266 3375 2271 3380
rect 2265 3314 2270 3319
rect 2443 3678 2447 3682
rect 2348 3518 2353 3523
rect 2323 3390 2328 3395
rect 2357 3383 2362 3388
rect 2354 3310 2359 3315
rect 1991 3190 1996 3195
rect 2027 3183 2032 3188
rect 2038 3187 2043 3192
rect 2061 3178 2066 3183
rect 2085 3183 2090 3188
rect 2114 3189 2119 3194
rect 2143 3189 2147 3194
rect 2100 3178 2105 3184
rect 2130 3183 2135 3188
rect 2159 3184 2164 3189
rect 2184 3178 2189 3183
rect 2241 3257 2246 3262
rect 2229 3189 2234 3194
rect 2288 3183 2293 3188
rect 2299 3187 2304 3192
rect 2322 3178 2327 3183
rect 2346 3183 2351 3188
rect 2375 3189 2380 3194
rect 2404 3189 2408 3194
rect 2361 3178 2366 3184
rect 2391 3183 2396 3188
rect 2416 3189 2421 3194
rect 2452 3190 2456 3194
rect 2290 3078 2294 3082
rect 2709 3693 2713 3697
rect 2415 2996 2419 3000
rect 1987 2747 1991 2751
rect 1989 2667 1994 2672
rect 2027 2664 2032 2669
rect 2038 2660 2043 2665
rect 2061 2669 2066 2674
rect 2085 2664 2090 2669
rect 2100 2668 2105 2674
rect 2130 2664 2135 2669
rect 2159 2663 2164 2668
rect 2114 2658 2119 2663
rect 2143 2658 2147 2663
rect 2185 2657 2190 2662
rect 1991 2604 1996 2609
rect 2027 2597 2032 2602
rect 2038 2601 2043 2606
rect 2061 2592 2066 2597
rect 2085 2597 2090 2602
rect 2114 2603 2119 2608
rect 2143 2603 2147 2608
rect 2100 2592 2105 2598
rect 2130 2597 2135 2602
rect 2159 2598 2164 2603
rect 2185 2598 2190 2603
rect 1990 2535 1995 2540
rect 2027 2532 2032 2537
rect 2038 2528 2043 2533
rect 2061 2537 2066 2542
rect 2085 2532 2090 2537
rect 2241 2663 2246 2668
rect 2100 2536 2105 2542
rect 2130 2532 2135 2537
rect 2159 2531 2164 2536
rect 2114 2526 2119 2531
rect 2143 2526 2147 2531
rect 2185 2525 2190 2530
rect 1991 2472 1996 2477
rect 2027 2465 2032 2470
rect 2038 2469 2043 2474
rect 2061 2460 2066 2465
rect 2085 2465 2090 2470
rect 2114 2471 2119 2476
rect 2143 2471 2147 2476
rect 2100 2460 2105 2466
rect 2130 2465 2135 2470
rect 2159 2466 2164 2471
rect 2184 2467 2189 2472
rect 1990 2403 1995 2408
rect 2027 2400 2032 2405
rect 2038 2396 2043 2401
rect 2061 2405 2066 2410
rect 2085 2400 2090 2405
rect 2100 2404 2105 2410
rect 2130 2400 2135 2405
rect 2159 2399 2164 2404
rect 2114 2394 2119 2399
rect 2143 2394 2147 2399
rect 2185 2393 2190 2398
rect 2241 2539 2246 2544
rect 2266 2657 2271 2662
rect 2265 2598 2270 2603
rect 2326 2663 2331 2668
rect 2290 2525 2295 2530
rect 2290 2467 2295 2472
rect 1991 2340 1996 2345
rect 2027 2333 2032 2338
rect 2038 2337 2043 2342
rect 2061 2328 2066 2333
rect 2085 2333 2090 2338
rect 2114 2339 2119 2344
rect 2143 2339 2147 2344
rect 2100 2328 2105 2334
rect 2130 2333 2135 2338
rect 2159 2334 2164 2339
rect 2185 2332 2190 2337
rect 1990 2271 1995 2276
rect 2027 2268 2032 2273
rect 2038 2264 2043 2269
rect 2061 2273 2066 2278
rect 2085 2268 2090 2273
rect 2100 2272 2105 2278
rect 2130 2268 2135 2273
rect 2159 2267 2164 2272
rect 2114 2262 2119 2267
rect 2143 2262 2147 2267
rect 2185 2261 2190 2266
rect 2241 2399 2246 2404
rect 2266 2393 2271 2398
rect 2265 2332 2270 2337
rect 2443 2696 2447 2700
rect 2708 3590 2712 3594
rect 2348 2536 2353 2541
rect 2323 2408 2328 2413
rect 2357 2401 2362 2406
rect 2354 2328 2359 2333
rect 1991 2208 1996 2213
rect 2027 2201 2032 2206
rect 2038 2205 2043 2210
rect 2061 2196 2066 2201
rect 2085 2201 2090 2206
rect 2114 2207 2119 2212
rect 2143 2207 2147 2212
rect 2100 2196 2105 2202
rect 2130 2201 2135 2206
rect 2159 2202 2164 2207
rect 2184 2196 2189 2201
rect 2241 2275 2246 2280
rect 2229 2207 2234 2212
rect 2288 2201 2293 2206
rect 2299 2205 2304 2210
rect 2322 2196 2327 2201
rect 2346 2201 2351 2206
rect 2375 2207 2380 2212
rect 2404 2207 2408 2212
rect 2361 2196 2366 2202
rect 2391 2201 2396 2206
rect 2416 2207 2421 2212
rect 2452 2208 2456 2212
rect 2290 2096 2294 2100
rect 2841 2823 2845 2827
rect 2709 2712 2713 2716
rect 2415 2014 2419 2018
rect 2708 2608 2712 2612
rect 2841 1841 2845 1845
rect 2932 3729 2936 3733
rect 2933 3649 2938 3654
rect 2972 3646 2977 3651
rect 2983 3642 2988 3647
rect 3006 3651 3011 3656
rect 3030 3646 3035 3651
rect 3045 3650 3050 3656
rect 3075 3646 3080 3651
rect 3104 3645 3109 3650
rect 3059 3640 3064 3645
rect 3088 3640 3092 3645
rect 3130 3639 3135 3644
rect 2936 3586 2941 3591
rect 2972 3579 2977 3584
rect 2983 3583 2988 3588
rect 3006 3574 3011 3579
rect 3030 3579 3035 3584
rect 3059 3585 3064 3590
rect 3088 3585 3092 3590
rect 3045 3574 3050 3580
rect 3075 3579 3080 3584
rect 3104 3580 3109 3585
rect 3130 3580 3135 3585
rect 2935 3517 2940 3522
rect 2972 3514 2977 3519
rect 2983 3510 2988 3515
rect 3006 3519 3011 3524
rect 3030 3514 3035 3519
rect 3186 3645 3191 3650
rect 3045 3518 3050 3524
rect 3075 3514 3080 3519
rect 3104 3513 3109 3518
rect 3059 3508 3064 3513
rect 3088 3508 3092 3513
rect 3130 3507 3135 3512
rect 2936 3454 2941 3459
rect 2972 3447 2977 3452
rect 2983 3451 2988 3456
rect 3006 3442 3011 3447
rect 3030 3447 3035 3452
rect 3059 3453 3064 3458
rect 3088 3453 3092 3458
rect 3045 3442 3050 3448
rect 3075 3447 3080 3452
rect 3104 3448 3109 3453
rect 3129 3449 3134 3454
rect 2935 3385 2940 3390
rect 2972 3382 2977 3387
rect 2983 3378 2988 3383
rect 3006 3387 3011 3392
rect 3030 3382 3035 3387
rect 3045 3386 3050 3392
rect 3075 3382 3080 3387
rect 3104 3381 3109 3386
rect 3059 3376 3064 3381
rect 3088 3376 3092 3381
rect 3130 3375 3135 3380
rect 3186 3521 3191 3526
rect 3211 3639 3216 3644
rect 3210 3580 3215 3585
rect 3271 3645 3276 3650
rect 3235 3507 3240 3512
rect 3235 3449 3240 3454
rect 2936 3322 2941 3327
rect 2972 3315 2977 3320
rect 2983 3319 2988 3324
rect 3006 3310 3011 3315
rect 3030 3315 3035 3320
rect 3059 3321 3064 3326
rect 3088 3321 3092 3326
rect 3045 3310 3050 3316
rect 3075 3315 3080 3320
rect 3104 3316 3109 3321
rect 3130 3314 3135 3319
rect 2935 3253 2940 3258
rect 2972 3250 2977 3255
rect 2983 3246 2988 3251
rect 3006 3255 3011 3260
rect 3030 3250 3035 3255
rect 3045 3254 3050 3260
rect 3075 3250 3080 3255
rect 3104 3249 3109 3254
rect 3059 3244 3064 3249
rect 3088 3244 3092 3249
rect 3130 3243 3135 3248
rect 3186 3381 3191 3386
rect 3211 3375 3216 3380
rect 3210 3314 3215 3319
rect 3388 3678 3392 3682
rect 3293 3518 3298 3523
rect 3268 3390 3273 3395
rect 3302 3383 3307 3388
rect 3299 3310 3304 3315
rect 2936 3190 2941 3195
rect 2972 3183 2977 3188
rect 2983 3187 2988 3192
rect 3006 3178 3011 3183
rect 3030 3183 3035 3188
rect 3059 3189 3064 3194
rect 3088 3189 3092 3194
rect 3045 3178 3050 3184
rect 3075 3183 3080 3188
rect 3104 3184 3109 3189
rect 3129 3178 3134 3183
rect 3186 3257 3191 3262
rect 3174 3189 3179 3194
rect 3233 3183 3238 3188
rect 3244 3187 3249 3192
rect 3267 3178 3272 3183
rect 3291 3183 3296 3188
rect 3320 3189 3325 3194
rect 3349 3189 3353 3194
rect 3306 3178 3311 3184
rect 3336 3183 3341 3188
rect 3361 3189 3366 3194
rect 3235 3078 3239 3082
rect 3360 2996 3364 3000
rect 2932 2747 2936 2751
rect 2934 2667 2939 2672
rect 2972 2664 2977 2669
rect 2983 2660 2988 2665
rect 3006 2669 3011 2674
rect 3030 2664 3035 2669
rect 3045 2668 3050 2674
rect 3075 2664 3080 2669
rect 3104 2663 3109 2668
rect 3059 2658 3064 2663
rect 3088 2658 3092 2663
rect 3130 2657 3135 2662
rect 2936 2604 2941 2609
rect 2972 2597 2977 2602
rect 2983 2601 2988 2606
rect 3006 2592 3011 2597
rect 3030 2597 3035 2602
rect 3059 2603 3064 2608
rect 3088 2603 3092 2608
rect 3045 2592 3050 2598
rect 3075 2597 3080 2602
rect 3104 2598 3109 2603
rect 3130 2598 3135 2603
rect 2935 2535 2940 2540
rect 2972 2532 2977 2537
rect 2983 2528 2988 2533
rect 3006 2537 3011 2542
rect 3030 2532 3035 2537
rect 3186 2663 3191 2668
rect 3045 2536 3050 2542
rect 3075 2532 3080 2537
rect 3104 2531 3109 2536
rect 3059 2526 3064 2531
rect 3088 2526 3092 2531
rect 3130 2525 3135 2530
rect 2936 2472 2941 2477
rect 2972 2465 2977 2470
rect 2983 2469 2988 2474
rect 3006 2460 3011 2465
rect 3030 2465 3035 2470
rect 3059 2471 3064 2476
rect 3088 2471 3092 2476
rect 3045 2460 3050 2466
rect 3075 2465 3080 2470
rect 3104 2466 3109 2471
rect 3129 2467 3134 2472
rect 2935 2403 2940 2408
rect 2972 2400 2977 2405
rect 2983 2396 2988 2401
rect 3006 2405 3011 2410
rect 3030 2400 3035 2405
rect 3045 2404 3050 2410
rect 3075 2400 3080 2405
rect 3104 2399 3109 2404
rect 3059 2394 3064 2399
rect 3088 2394 3092 2399
rect 3130 2393 3135 2398
rect 3186 2539 3191 2544
rect 3211 2657 3216 2662
rect 3210 2598 3215 2603
rect 3271 2663 3276 2668
rect 3235 2525 3240 2530
rect 3235 2467 3240 2472
rect 2936 2340 2941 2345
rect 2972 2333 2977 2338
rect 2983 2337 2988 2342
rect 3006 2328 3011 2333
rect 3030 2333 3035 2338
rect 3059 2339 3064 2344
rect 3088 2339 3092 2344
rect 3045 2328 3050 2334
rect 3075 2333 3080 2338
rect 3104 2334 3109 2339
rect 3130 2332 3135 2337
rect 2935 2271 2940 2276
rect 2972 2268 2977 2273
rect 2983 2264 2988 2269
rect 3006 2273 3011 2278
rect 3030 2268 3035 2273
rect 3045 2272 3050 2278
rect 3075 2268 3080 2273
rect 3104 2267 3109 2272
rect 3059 2262 3064 2267
rect 3088 2262 3092 2267
rect 3130 2261 3135 2266
rect 3186 2399 3191 2404
rect 3211 2393 3216 2398
rect 3210 2332 3215 2337
rect 3388 2696 3392 2700
rect 3293 2536 3298 2541
rect 3268 2408 3273 2413
rect 3302 2401 3307 2406
rect 3299 2328 3304 2333
rect 2936 2208 2941 2213
rect 2972 2201 2977 2206
rect 2983 2205 2988 2210
rect 3006 2196 3011 2201
rect 3030 2201 3035 2206
rect 3059 2207 3064 2212
rect 3088 2207 3092 2212
rect 3045 2196 3050 2202
rect 3075 2201 3080 2206
rect 3104 2202 3109 2207
rect 3129 2196 3134 2201
rect 3186 2275 3191 2280
rect 3174 2207 3179 2212
rect 3233 2201 3238 2206
rect 3244 2205 3249 2210
rect 3267 2196 3272 2201
rect 3291 2201 3296 2206
rect 3320 2207 3325 2212
rect 3349 2207 3353 2212
rect 3306 2196 3311 2202
rect 3336 2201 3341 2206
rect 3361 2207 3366 2212
rect 3235 2096 3239 2100
rect 3360 2014 3364 2018
<< metal3 >>
rect 2080 4448 2088 4450
rect 2080 4443 2081 4448
rect 2086 4443 2088 4448
rect 2080 4442 2088 4443
rect 2171 4330 2177 4331
rect 2171 4326 2172 4330
rect 2176 4326 2177 4330
rect 2171 4325 2177 4326
rect 1986 3733 1992 3734
rect 1986 3729 1987 3733
rect 1991 3729 1992 3733
rect 1986 3728 1992 3729
rect 2931 3733 2937 3734
rect 2931 3729 2932 3733
rect 2936 3729 2937 3733
rect 2931 3728 2937 3729
rect 1986 3698 1991 3728
rect 2931 3698 2936 3728
rect 1763 3697 1991 3698
rect 1763 3693 1764 3697
rect 1768 3693 1991 3697
rect 2708 3697 2936 3698
rect 2708 3693 2709 3697
rect 2713 3693 2936 3697
rect 1763 3692 1769 3693
rect 2708 3692 2714 3693
rect 2442 3682 2448 3683
rect 2442 3678 2443 3682
rect 2447 3678 2448 3682
rect 2442 3677 2448 3678
rect 3387 3682 3393 3683
rect 3387 3678 3388 3682
rect 3392 3678 3393 3682
rect 3387 3677 3393 3678
rect 2027 3656 2067 3657
rect 2027 3652 2061 3656
rect 2026 3651 2033 3652
rect 2026 3646 2027 3651
rect 2032 3646 2033 3651
rect 2060 3651 2061 3652
rect 2066 3651 2067 3656
rect 2099 3656 2135 3661
rect 2060 3650 2067 3651
rect 2084 3651 2091 3652
rect 2026 3645 2033 3646
rect 2037 3647 2044 3648
rect 2037 3642 2038 3647
rect 2043 3642 2044 3647
rect 2084 3646 2085 3651
rect 2090 3646 2091 3651
rect 2099 3650 2100 3656
rect 2105 3655 2135 3656
rect 2105 3650 2106 3655
rect 2130 3652 2135 3655
rect 2099 3649 2106 3650
rect 2129 3651 2136 3652
rect 2129 3646 2130 3651
rect 2135 3646 2136 3651
rect 2158 3650 2165 3651
rect 2084 3645 2091 3646
rect 2113 3645 2120 3646
rect 2129 3645 2136 3646
rect 2142 3645 2148 3646
rect 2085 3642 2090 3645
rect 2037 3637 2090 3642
rect 2113 3640 2114 3645
rect 2119 3640 2120 3645
rect 2142 3640 2143 3645
rect 2147 3640 2148 3645
rect 2113 3639 2148 3640
rect 2114 3635 2148 3639
rect 2158 3645 2159 3650
rect 2164 3645 2165 3650
rect 2240 3650 2247 3651
rect 2240 3645 2241 3650
rect 2246 3645 2247 3650
rect 2325 3650 2332 3651
rect 2325 3645 2326 3650
rect 2331 3645 2332 3650
rect 2158 3644 2165 3645
rect 2184 3644 2191 3645
rect 2240 3644 2247 3645
rect 2265 3644 2272 3645
rect 2325 3644 2332 3645
rect 2158 3639 2185 3644
rect 2190 3639 2191 3644
rect 2241 3639 2266 3644
rect 2271 3639 2272 3644
rect 2158 3618 2163 3639
rect 2184 3638 2191 3639
rect 2265 3638 2272 3639
rect 2322 3639 2331 3644
rect 1991 3612 2163 3618
rect 1762 3594 1768 3595
rect 1762 3590 1763 3594
rect 1767 3590 1900 3594
rect 1991 3592 1996 3612
rect 1762 3589 1900 3590
rect 1506 3194 1512 3195
rect 1506 3190 1507 3194
rect 1511 3190 1512 3194
rect 1506 3189 1512 3190
rect 1895 2828 1900 3589
rect 1990 3591 1997 3592
rect 1990 3586 1991 3591
rect 1996 3586 1997 3591
rect 1990 3585 1997 3586
rect 2037 3588 2090 3593
rect 2114 3591 2148 3595
rect 2026 3584 2033 3585
rect 2026 3579 2027 3584
rect 2032 3579 2033 3584
rect 2037 3583 2038 3588
rect 2043 3583 2044 3588
rect 2085 3585 2090 3588
rect 2113 3590 2148 3591
rect 2113 3585 2114 3590
rect 2119 3585 2120 3590
rect 2142 3585 2143 3590
rect 2147 3585 2148 3590
rect 2037 3582 2044 3583
rect 2084 3584 2091 3585
rect 2113 3584 2120 3585
rect 2129 3584 2136 3585
rect 2142 3584 2148 3585
rect 2158 3585 2165 3586
rect 2184 3585 2191 3586
rect 2264 3585 2271 3586
rect 2026 3578 2033 3579
rect 2060 3579 2067 3580
rect 2060 3578 2061 3579
rect 2027 3574 2061 3578
rect 2066 3574 2067 3579
rect 2084 3579 2085 3584
rect 2090 3579 2091 3584
rect 2084 3578 2091 3579
rect 2099 3580 2106 3581
rect 2027 3573 2067 3574
rect 2099 3574 2100 3580
rect 2105 3575 2106 3580
rect 2129 3579 2130 3584
rect 2135 3579 2136 3584
rect 2158 3580 2159 3585
rect 2164 3580 2185 3585
rect 2190 3580 2191 3585
rect 2158 3579 2165 3580
rect 2184 3579 2191 3580
rect 2241 3580 2265 3585
rect 2270 3580 2271 3585
rect 2129 3578 2136 3579
rect 2130 3575 2135 3578
rect 2105 3574 2135 3575
rect 2099 3569 2135 3574
rect 2159 3552 2164 3579
rect 1990 3546 2164 3552
rect 1990 3523 1995 3546
rect 2027 3524 2067 3525
rect 1989 3522 1996 3523
rect 1989 3517 1990 3522
rect 1995 3517 1996 3522
rect 2027 3520 2061 3524
rect 1989 3516 1996 3517
rect 2026 3519 2033 3520
rect 2026 3514 2027 3519
rect 2032 3514 2033 3519
rect 2060 3519 2061 3520
rect 2066 3519 2067 3524
rect 2099 3524 2135 3529
rect 2241 3527 2246 3580
rect 2264 3579 2271 3580
rect 2322 3551 2327 3639
rect 2284 3546 2327 3551
rect 2060 3518 2067 3519
rect 2084 3519 2091 3520
rect 2026 3513 2033 3514
rect 2037 3515 2044 3516
rect 2037 3510 2038 3515
rect 2043 3510 2044 3515
rect 2084 3514 2085 3519
rect 2090 3514 2091 3519
rect 2099 3518 2100 3524
rect 2105 3523 2135 3524
rect 2105 3518 2106 3523
rect 2130 3520 2135 3523
rect 2240 3526 2247 3527
rect 2240 3521 2241 3526
rect 2246 3521 2247 3526
rect 2240 3520 2247 3521
rect 2099 3517 2106 3518
rect 2129 3519 2136 3520
rect 2129 3514 2130 3519
rect 2135 3514 2136 3519
rect 2158 3518 2165 3519
rect 2084 3513 2091 3514
rect 2113 3513 2120 3514
rect 2129 3513 2136 3514
rect 2142 3513 2148 3514
rect 2085 3510 2090 3513
rect 2037 3505 2090 3510
rect 2113 3508 2114 3513
rect 2119 3508 2120 3513
rect 2142 3508 2143 3513
rect 2147 3508 2148 3513
rect 2113 3507 2148 3508
rect 2114 3503 2148 3507
rect 2158 3513 2159 3518
rect 2164 3513 2165 3518
rect 2284 3513 2289 3546
rect 2347 3523 2354 3524
rect 2347 3518 2348 3523
rect 2353 3518 2354 3523
rect 2347 3517 2354 3518
rect 2158 3512 2165 3513
rect 2184 3512 2191 3513
rect 2158 3507 2185 3512
rect 2190 3507 2191 3512
rect 2284 3512 2296 3513
rect 2284 3507 2290 3512
rect 2295 3507 2296 3512
rect 2158 3486 2163 3507
rect 2184 3506 2191 3507
rect 2289 3506 2296 3507
rect 1991 3480 2163 3486
rect 1991 3460 1996 3480
rect 1990 3459 1997 3460
rect 1990 3454 1991 3459
rect 1996 3454 1997 3459
rect 1990 3453 1997 3454
rect 2037 3456 2090 3461
rect 2114 3459 2148 3463
rect 2026 3452 2033 3453
rect 2026 3447 2027 3452
rect 2032 3447 2033 3452
rect 2037 3451 2038 3456
rect 2043 3451 2044 3456
rect 2085 3453 2090 3456
rect 2113 3458 2148 3459
rect 2113 3453 2114 3458
rect 2119 3453 2120 3458
rect 2142 3453 2143 3458
rect 2147 3453 2148 3458
rect 2183 3454 2190 3455
rect 2289 3454 2296 3455
rect 2037 3450 2044 3451
rect 2084 3452 2091 3453
rect 2113 3452 2120 3453
rect 2129 3452 2136 3453
rect 2142 3452 2148 3453
rect 2158 3453 2184 3454
rect 2026 3446 2033 3447
rect 2060 3447 2067 3448
rect 2060 3446 2061 3447
rect 2027 3442 2061 3446
rect 2066 3442 2067 3447
rect 2084 3447 2085 3452
rect 2090 3447 2091 3452
rect 2084 3446 2091 3447
rect 2099 3448 2106 3449
rect 2027 3441 2067 3442
rect 2099 3442 2100 3448
rect 2105 3443 2106 3448
rect 2129 3447 2130 3452
rect 2135 3447 2136 3452
rect 2129 3446 2136 3447
rect 2158 3448 2159 3453
rect 2164 3449 2184 3453
rect 2189 3449 2190 3454
rect 2164 3448 2165 3449
rect 2183 3448 2190 3449
rect 2285 3449 2290 3454
rect 2295 3449 2296 3454
rect 2285 3448 2296 3449
rect 2158 3447 2165 3448
rect 2130 3443 2135 3446
rect 2105 3442 2135 3443
rect 2099 3437 2135 3442
rect 2158 3420 2163 3447
rect 1990 3414 2163 3420
rect 2285 3420 2290 3448
rect 2285 3415 2328 3420
rect 1990 3391 1995 3414
rect 2027 3392 2067 3393
rect 1989 3390 1996 3391
rect 1989 3385 1990 3390
rect 1995 3385 1996 3390
rect 2027 3388 2061 3392
rect 1989 3384 1996 3385
rect 2026 3387 2033 3388
rect 2026 3382 2027 3387
rect 2032 3382 2033 3387
rect 2060 3387 2061 3388
rect 2066 3387 2067 3392
rect 2099 3392 2135 3397
rect 2323 3396 2328 3415
rect 2060 3386 2067 3387
rect 2084 3387 2091 3388
rect 2026 3381 2033 3382
rect 2037 3383 2044 3384
rect 2037 3378 2038 3383
rect 2043 3378 2044 3383
rect 2084 3382 2085 3387
rect 2090 3382 2091 3387
rect 2099 3386 2100 3392
rect 2105 3391 2135 3392
rect 2105 3386 2106 3391
rect 2130 3388 2135 3391
rect 2322 3395 2329 3396
rect 2322 3390 2323 3395
rect 2328 3390 2329 3395
rect 2322 3389 2329 3390
rect 2348 3388 2353 3517
rect 2356 3388 2363 3389
rect 2099 3385 2106 3386
rect 2129 3387 2136 3388
rect 2129 3382 2130 3387
rect 2135 3382 2136 3387
rect 2158 3386 2165 3387
rect 2084 3381 2091 3382
rect 2113 3381 2120 3382
rect 2129 3381 2136 3382
rect 2142 3381 2148 3382
rect 2085 3378 2090 3381
rect 2037 3373 2090 3378
rect 2113 3376 2114 3381
rect 2119 3376 2120 3381
rect 2142 3376 2143 3381
rect 2147 3376 2148 3381
rect 2113 3375 2148 3376
rect 2114 3371 2148 3375
rect 2158 3381 2159 3386
rect 2164 3381 2165 3386
rect 2240 3386 2247 3387
rect 2240 3381 2241 3386
rect 2246 3381 2247 3386
rect 2336 3383 2357 3388
rect 2362 3383 2363 3388
rect 2336 3382 2348 3383
rect 2356 3382 2363 3383
rect 2158 3380 2165 3381
rect 2184 3380 2191 3381
rect 2240 3380 2247 3381
rect 2265 3380 2272 3381
rect 2158 3375 2185 3380
rect 2190 3375 2191 3380
rect 2241 3375 2266 3380
rect 2271 3375 2272 3380
rect 2158 3354 2163 3375
rect 2184 3374 2191 3375
rect 2265 3374 2272 3375
rect 2336 3374 2341 3382
rect 1991 3348 2163 3354
rect 2303 3353 2341 3374
rect 1991 3328 1996 3348
rect 1990 3327 1997 3328
rect 1990 3322 1991 3327
rect 1996 3322 1997 3327
rect 1990 3321 1997 3322
rect 2037 3324 2090 3329
rect 2114 3327 2148 3331
rect 2026 3320 2033 3321
rect 2026 3315 2027 3320
rect 2032 3315 2033 3320
rect 2037 3319 2038 3324
rect 2043 3319 2044 3324
rect 2085 3321 2090 3324
rect 2113 3326 2148 3327
rect 2113 3321 2114 3326
rect 2119 3321 2120 3326
rect 2142 3321 2143 3326
rect 2147 3321 2148 3326
rect 2037 3318 2044 3319
rect 2084 3320 2091 3321
rect 2113 3320 2120 3321
rect 2129 3320 2136 3321
rect 2142 3320 2148 3321
rect 2158 3321 2165 3322
rect 2026 3314 2033 3315
rect 2060 3315 2067 3316
rect 2060 3314 2061 3315
rect 2027 3310 2061 3314
rect 2066 3310 2067 3315
rect 2084 3315 2085 3320
rect 2090 3315 2091 3320
rect 2084 3314 2091 3315
rect 2099 3316 2106 3317
rect 2027 3309 2067 3310
rect 2099 3310 2100 3316
rect 2105 3311 2106 3316
rect 2129 3315 2130 3320
rect 2135 3315 2136 3320
rect 2158 3316 2159 3321
rect 2164 3319 2165 3321
rect 2184 3319 2191 3320
rect 2264 3319 2271 3320
rect 2164 3316 2185 3319
rect 2158 3315 2185 3316
rect 2129 3314 2136 3315
rect 2159 3314 2185 3315
rect 2190 3314 2191 3319
rect 2130 3311 2135 3314
rect 2105 3310 2135 3311
rect 2099 3305 2135 3310
rect 2159 3288 2164 3314
rect 2184 3313 2191 3314
rect 2241 3314 2265 3319
rect 2270 3314 2271 3319
rect 1990 3282 2164 3288
rect 1990 3259 1995 3282
rect 2027 3260 2067 3261
rect 1989 3258 1996 3259
rect 1989 3253 1990 3258
rect 1995 3253 1996 3258
rect 2027 3256 2061 3260
rect 1989 3252 1996 3253
rect 2026 3255 2033 3256
rect 2026 3250 2027 3255
rect 2032 3250 2033 3255
rect 2060 3255 2061 3256
rect 2066 3255 2067 3260
rect 2099 3260 2135 3265
rect 2241 3263 2246 3314
rect 2264 3313 2271 3314
rect 2060 3254 2067 3255
rect 2084 3255 2091 3256
rect 2026 3249 2033 3250
rect 2037 3251 2044 3252
rect 2037 3246 2038 3251
rect 2043 3246 2044 3251
rect 2084 3250 2085 3255
rect 2090 3250 2091 3255
rect 2099 3254 2100 3260
rect 2105 3259 2135 3260
rect 2105 3254 2106 3259
rect 2130 3256 2135 3259
rect 2240 3262 2247 3263
rect 2240 3257 2241 3262
rect 2246 3257 2247 3262
rect 2240 3256 2247 3257
rect 2099 3253 2106 3254
rect 2129 3255 2136 3256
rect 2129 3250 2130 3255
rect 2135 3250 2136 3255
rect 2158 3254 2165 3255
rect 2084 3249 2091 3250
rect 2113 3249 2120 3250
rect 2129 3249 2136 3250
rect 2142 3249 2148 3250
rect 2085 3246 2090 3249
rect 2037 3241 2090 3246
rect 2113 3244 2114 3249
rect 2119 3244 2120 3249
rect 2142 3244 2143 3249
rect 2147 3244 2148 3249
rect 2113 3243 2148 3244
rect 2114 3239 2148 3243
rect 2158 3249 2159 3254
rect 2164 3249 2165 3254
rect 2158 3248 2165 3249
rect 2184 3248 2191 3249
rect 2158 3243 2185 3248
rect 2190 3243 2191 3248
rect 2303 3244 2308 3353
rect 2353 3315 2360 3316
rect 2353 3310 2354 3315
rect 2359 3310 2360 3315
rect 2353 3309 2360 3310
rect 2260 3243 2308 3244
rect 2158 3222 2163 3243
rect 2184 3242 2191 3243
rect 1991 3216 2163 3222
rect 2229 3238 2308 3243
rect 2354 3247 2359 3309
rect 2354 3241 2421 3247
rect 1991 3196 1996 3216
rect 1990 3195 1997 3196
rect 1990 3190 1991 3195
rect 1996 3190 1997 3195
rect 1990 3189 1997 3190
rect 2037 3192 2090 3197
rect 2114 3195 2148 3199
rect 2229 3195 2234 3238
rect 2026 3188 2033 3189
rect 2026 3183 2027 3188
rect 2032 3183 2033 3188
rect 2037 3187 2038 3192
rect 2043 3187 2044 3192
rect 2085 3189 2090 3192
rect 2113 3194 2148 3195
rect 2113 3189 2114 3194
rect 2119 3189 2120 3194
rect 2142 3189 2143 3194
rect 2147 3189 2148 3194
rect 2228 3194 2235 3195
rect 2037 3186 2044 3187
rect 2084 3188 2091 3189
rect 2113 3188 2120 3189
rect 2129 3188 2136 3189
rect 2142 3188 2148 3189
rect 2158 3189 2165 3190
rect 2026 3182 2033 3183
rect 2060 3183 2067 3184
rect 2060 3182 2061 3183
rect 2027 3178 2061 3182
rect 2066 3178 2067 3183
rect 2084 3183 2085 3188
rect 2090 3183 2091 3188
rect 2084 3182 2091 3183
rect 2099 3184 2106 3185
rect 2027 3177 2067 3178
rect 2099 3178 2100 3184
rect 2105 3179 2106 3184
rect 2129 3183 2130 3188
rect 2135 3183 2136 3188
rect 2158 3184 2159 3189
rect 2164 3184 2165 3189
rect 2228 3189 2229 3194
rect 2234 3189 2235 3194
rect 2298 3192 2351 3197
rect 2375 3195 2409 3199
rect 2416 3195 2421 3241
rect 2228 3188 2235 3189
rect 2287 3188 2294 3189
rect 2158 3183 2165 3184
rect 2183 3183 2190 3184
rect 2129 3182 2136 3183
rect 2130 3179 2135 3182
rect 2105 3178 2135 3179
rect 2099 3173 2135 3178
rect 2160 3178 2184 3183
rect 2189 3178 2190 3183
rect 2287 3183 2288 3188
rect 2293 3183 2294 3188
rect 2298 3187 2299 3192
rect 2304 3187 2305 3192
rect 2346 3189 2351 3192
rect 2374 3194 2409 3195
rect 2374 3189 2375 3194
rect 2380 3189 2381 3194
rect 2403 3189 2404 3194
rect 2408 3189 2409 3194
rect 2298 3186 2305 3187
rect 2345 3188 2352 3189
rect 2374 3188 2381 3189
rect 2390 3188 2397 3189
rect 2403 3188 2409 3189
rect 2415 3194 2422 3195
rect 2415 3189 2416 3194
rect 2421 3189 2422 3194
rect 2415 3188 2422 3189
rect 2287 3182 2294 3183
rect 2321 3183 2328 3184
rect 2321 3182 2322 3183
rect 1895 2827 1901 2828
rect 1895 2823 1896 2827
rect 1900 2823 1901 2827
rect 1895 2822 1901 2823
rect 2160 2810 2165 3178
rect 2183 3177 2190 3178
rect 2288 3178 2322 3182
rect 2327 3178 2328 3183
rect 2345 3183 2346 3188
rect 2351 3183 2352 3188
rect 2345 3182 2352 3183
rect 2360 3184 2367 3185
rect 2288 3177 2328 3178
rect 2360 3178 2361 3184
rect 2366 3179 2367 3184
rect 2390 3183 2391 3188
rect 2396 3183 2397 3188
rect 2390 3182 2397 3183
rect 2391 3179 2396 3182
rect 2366 3178 2396 3179
rect 2360 3173 2396 3178
rect 2443 3150 2448 3677
rect 2972 3656 3012 3657
rect 2932 3654 2939 3655
rect 2910 3649 2933 3654
rect 2938 3649 2939 3654
rect 2972 3652 3006 3656
rect 2707 3594 2713 3595
rect 2707 3590 2708 3594
rect 2712 3590 2845 3594
rect 2707 3589 2845 3590
rect 2451 3194 2457 3195
rect 2451 3190 2452 3194
rect 2456 3190 2457 3194
rect 2451 3189 2457 3190
rect 2290 3145 2448 3150
rect 2290 3083 2295 3145
rect 2289 3082 2295 3083
rect 2289 3078 2290 3082
rect 2294 3078 2295 3082
rect 2289 3077 2295 3078
rect 2452 3020 2457 3189
rect 2415 3015 2457 3020
rect 2415 3001 2420 3015
rect 2414 3000 2420 3001
rect 2414 2996 2415 3000
rect 2419 2996 2420 3000
rect 2414 2995 2420 2996
rect 2840 2828 2845 3589
rect 2840 2827 2846 2828
rect 2840 2823 2841 2827
rect 2845 2823 2846 2827
rect 2840 2822 2846 2823
rect 2910 2810 2915 3649
rect 2932 3648 2939 3649
rect 2971 3651 2978 3652
rect 2971 3646 2972 3651
rect 2977 3646 2978 3651
rect 3005 3651 3006 3652
rect 3011 3651 3012 3656
rect 3044 3656 3080 3661
rect 3005 3650 3012 3651
rect 3029 3651 3036 3652
rect 2971 3645 2978 3646
rect 2982 3647 2989 3648
rect 2982 3642 2983 3647
rect 2988 3642 2989 3647
rect 3029 3646 3030 3651
rect 3035 3646 3036 3651
rect 3044 3650 3045 3656
rect 3050 3655 3080 3656
rect 3050 3650 3051 3655
rect 3075 3652 3080 3655
rect 3044 3649 3051 3650
rect 3074 3651 3081 3652
rect 3074 3646 3075 3651
rect 3080 3646 3081 3651
rect 3103 3650 3110 3651
rect 3029 3645 3036 3646
rect 3058 3645 3065 3646
rect 3074 3645 3081 3646
rect 3087 3645 3093 3646
rect 3030 3642 3035 3645
rect 2982 3637 3035 3642
rect 3058 3640 3059 3645
rect 3064 3640 3065 3645
rect 3087 3640 3088 3645
rect 3092 3640 3093 3645
rect 3058 3639 3093 3640
rect 3059 3635 3093 3639
rect 3103 3645 3104 3650
rect 3109 3645 3110 3650
rect 3185 3650 3192 3651
rect 3185 3645 3186 3650
rect 3191 3645 3192 3650
rect 3270 3650 3277 3651
rect 3270 3645 3271 3650
rect 3276 3645 3277 3650
rect 3103 3644 3110 3645
rect 3129 3644 3136 3645
rect 3185 3644 3192 3645
rect 3210 3644 3217 3645
rect 3270 3644 3277 3645
rect 3103 3639 3130 3644
rect 3135 3639 3136 3644
rect 3186 3639 3211 3644
rect 3216 3639 3217 3644
rect 3103 3618 3108 3639
rect 3129 3638 3136 3639
rect 3210 3638 3217 3639
rect 3267 3639 3276 3644
rect 2936 3612 3108 3618
rect 2936 3592 2941 3612
rect 2935 3591 2942 3592
rect 2935 3586 2936 3591
rect 2941 3586 2942 3591
rect 2935 3585 2942 3586
rect 2982 3588 3035 3593
rect 3059 3591 3093 3595
rect 2971 3584 2978 3585
rect 2971 3579 2972 3584
rect 2977 3579 2978 3584
rect 2982 3583 2983 3588
rect 2988 3583 2989 3588
rect 3030 3585 3035 3588
rect 3058 3590 3093 3591
rect 3058 3585 3059 3590
rect 3064 3585 3065 3590
rect 3087 3585 3088 3590
rect 3092 3585 3093 3590
rect 2982 3582 2989 3583
rect 3029 3584 3036 3585
rect 3058 3584 3065 3585
rect 3074 3584 3081 3585
rect 3087 3584 3093 3585
rect 3103 3585 3110 3586
rect 3129 3585 3136 3586
rect 3209 3585 3216 3586
rect 2971 3578 2978 3579
rect 3005 3579 3012 3580
rect 3005 3578 3006 3579
rect 2972 3574 3006 3578
rect 3011 3574 3012 3579
rect 3029 3579 3030 3584
rect 3035 3579 3036 3584
rect 3029 3578 3036 3579
rect 3044 3580 3051 3581
rect 2972 3573 3012 3574
rect 3044 3574 3045 3580
rect 3050 3575 3051 3580
rect 3074 3579 3075 3584
rect 3080 3579 3081 3584
rect 3103 3580 3104 3585
rect 3109 3580 3130 3585
rect 3135 3580 3136 3585
rect 3103 3579 3110 3580
rect 3129 3579 3136 3580
rect 3186 3580 3210 3585
rect 3215 3580 3216 3585
rect 3074 3578 3081 3579
rect 3075 3575 3080 3578
rect 3050 3574 3080 3575
rect 3044 3569 3080 3574
rect 3104 3552 3109 3579
rect 2935 3546 3109 3552
rect 2935 3523 2940 3546
rect 2972 3524 3012 3525
rect 2934 3522 2941 3523
rect 2934 3517 2935 3522
rect 2940 3517 2941 3522
rect 2972 3520 3006 3524
rect 2934 3516 2941 3517
rect 2971 3519 2978 3520
rect 2971 3514 2972 3519
rect 2977 3514 2978 3519
rect 3005 3519 3006 3520
rect 3011 3519 3012 3524
rect 3044 3524 3080 3529
rect 3186 3527 3191 3580
rect 3209 3579 3216 3580
rect 3267 3551 3272 3639
rect 3229 3546 3272 3551
rect 3005 3518 3012 3519
rect 3029 3519 3036 3520
rect 2971 3513 2978 3514
rect 2982 3515 2989 3516
rect 2982 3510 2983 3515
rect 2988 3510 2989 3515
rect 3029 3514 3030 3519
rect 3035 3514 3036 3519
rect 3044 3518 3045 3524
rect 3050 3523 3080 3524
rect 3050 3518 3051 3523
rect 3075 3520 3080 3523
rect 3185 3526 3192 3527
rect 3185 3521 3186 3526
rect 3191 3521 3192 3526
rect 3185 3520 3192 3521
rect 3044 3517 3051 3518
rect 3074 3519 3081 3520
rect 3074 3514 3075 3519
rect 3080 3514 3081 3519
rect 3103 3518 3110 3519
rect 3029 3513 3036 3514
rect 3058 3513 3065 3514
rect 3074 3513 3081 3514
rect 3087 3513 3093 3514
rect 3030 3510 3035 3513
rect 2982 3505 3035 3510
rect 3058 3508 3059 3513
rect 3064 3508 3065 3513
rect 3087 3508 3088 3513
rect 3092 3508 3093 3513
rect 3058 3507 3093 3508
rect 3059 3503 3093 3507
rect 3103 3513 3104 3518
rect 3109 3513 3110 3518
rect 3229 3513 3234 3546
rect 3292 3523 3299 3524
rect 3292 3518 3293 3523
rect 3298 3518 3299 3523
rect 3292 3517 3299 3518
rect 3103 3512 3110 3513
rect 3129 3512 3136 3513
rect 3103 3507 3130 3512
rect 3135 3507 3136 3512
rect 3229 3512 3241 3513
rect 3229 3507 3235 3512
rect 3240 3507 3241 3512
rect 3103 3486 3108 3507
rect 3129 3506 3136 3507
rect 3234 3506 3241 3507
rect 2936 3480 3108 3486
rect 2936 3460 2941 3480
rect 2935 3459 2942 3460
rect 2935 3454 2936 3459
rect 2941 3454 2942 3459
rect 2935 3453 2942 3454
rect 2982 3456 3035 3461
rect 3059 3459 3093 3463
rect 2971 3452 2978 3453
rect 2971 3447 2972 3452
rect 2977 3447 2978 3452
rect 2982 3451 2983 3456
rect 2988 3451 2989 3456
rect 3030 3453 3035 3456
rect 3058 3458 3093 3459
rect 3058 3453 3059 3458
rect 3064 3453 3065 3458
rect 3087 3453 3088 3458
rect 3092 3453 3093 3458
rect 3128 3454 3135 3455
rect 3234 3454 3241 3455
rect 2982 3450 2989 3451
rect 3029 3452 3036 3453
rect 3058 3452 3065 3453
rect 3074 3452 3081 3453
rect 3087 3452 3093 3453
rect 3103 3453 3129 3454
rect 2971 3446 2978 3447
rect 3005 3447 3012 3448
rect 3005 3446 3006 3447
rect 2972 3442 3006 3446
rect 3011 3442 3012 3447
rect 3029 3447 3030 3452
rect 3035 3447 3036 3452
rect 3029 3446 3036 3447
rect 3044 3448 3051 3449
rect 2972 3441 3012 3442
rect 3044 3442 3045 3448
rect 3050 3443 3051 3448
rect 3074 3447 3075 3452
rect 3080 3447 3081 3452
rect 3074 3446 3081 3447
rect 3103 3448 3104 3453
rect 3109 3449 3129 3453
rect 3134 3449 3135 3454
rect 3109 3448 3110 3449
rect 3128 3448 3135 3449
rect 3230 3449 3235 3454
rect 3240 3449 3241 3454
rect 3230 3448 3241 3449
rect 3103 3447 3110 3448
rect 3075 3443 3080 3446
rect 3050 3442 3080 3443
rect 3044 3437 3080 3442
rect 3103 3420 3108 3447
rect 2935 3414 3108 3420
rect 3230 3420 3235 3448
rect 3230 3415 3273 3420
rect 2935 3391 2940 3414
rect 2972 3392 3012 3393
rect 2934 3390 2941 3391
rect 2934 3385 2935 3390
rect 2940 3385 2941 3390
rect 2972 3388 3006 3392
rect 2934 3384 2941 3385
rect 2971 3387 2978 3388
rect 2971 3382 2972 3387
rect 2977 3382 2978 3387
rect 3005 3387 3006 3388
rect 3011 3387 3012 3392
rect 3044 3392 3080 3397
rect 3268 3396 3273 3415
rect 3005 3386 3012 3387
rect 3029 3387 3036 3388
rect 2971 3381 2978 3382
rect 2982 3383 2989 3384
rect 2982 3378 2983 3383
rect 2988 3378 2989 3383
rect 3029 3382 3030 3387
rect 3035 3382 3036 3387
rect 3044 3386 3045 3392
rect 3050 3391 3080 3392
rect 3050 3386 3051 3391
rect 3075 3388 3080 3391
rect 3267 3395 3274 3396
rect 3267 3390 3268 3395
rect 3273 3390 3274 3395
rect 3267 3389 3274 3390
rect 3293 3388 3298 3517
rect 3301 3388 3308 3389
rect 3044 3385 3051 3386
rect 3074 3387 3081 3388
rect 3074 3382 3075 3387
rect 3080 3382 3081 3387
rect 3103 3386 3110 3387
rect 3029 3381 3036 3382
rect 3058 3381 3065 3382
rect 3074 3381 3081 3382
rect 3087 3381 3093 3382
rect 3030 3378 3035 3381
rect 2982 3373 3035 3378
rect 3058 3376 3059 3381
rect 3064 3376 3065 3381
rect 3087 3376 3088 3381
rect 3092 3376 3093 3381
rect 3058 3375 3093 3376
rect 3059 3371 3093 3375
rect 3103 3381 3104 3386
rect 3109 3381 3110 3386
rect 3185 3386 3192 3387
rect 3185 3381 3186 3386
rect 3191 3381 3192 3386
rect 3281 3383 3302 3388
rect 3307 3383 3308 3388
rect 3281 3382 3293 3383
rect 3301 3382 3308 3383
rect 3103 3380 3110 3381
rect 3129 3380 3136 3381
rect 3185 3380 3192 3381
rect 3210 3380 3217 3381
rect 3103 3375 3130 3380
rect 3135 3375 3136 3380
rect 3186 3375 3211 3380
rect 3216 3375 3217 3380
rect 3103 3354 3108 3375
rect 3129 3374 3136 3375
rect 3210 3374 3217 3375
rect 3281 3374 3286 3382
rect 2936 3348 3108 3354
rect 3248 3353 3286 3374
rect 2936 3328 2941 3348
rect 2935 3327 2942 3328
rect 2935 3322 2936 3327
rect 2941 3322 2942 3327
rect 2935 3321 2942 3322
rect 2982 3324 3035 3329
rect 3059 3327 3093 3331
rect 2971 3320 2978 3321
rect 2971 3315 2972 3320
rect 2977 3315 2978 3320
rect 2982 3319 2983 3324
rect 2988 3319 2989 3324
rect 3030 3321 3035 3324
rect 3058 3326 3093 3327
rect 3058 3321 3059 3326
rect 3064 3321 3065 3326
rect 3087 3321 3088 3326
rect 3092 3321 3093 3326
rect 2982 3318 2989 3319
rect 3029 3320 3036 3321
rect 3058 3320 3065 3321
rect 3074 3320 3081 3321
rect 3087 3320 3093 3321
rect 3103 3321 3110 3322
rect 2971 3314 2978 3315
rect 3005 3315 3012 3316
rect 3005 3314 3006 3315
rect 2972 3310 3006 3314
rect 3011 3310 3012 3315
rect 3029 3315 3030 3320
rect 3035 3315 3036 3320
rect 3029 3314 3036 3315
rect 3044 3316 3051 3317
rect 2972 3309 3012 3310
rect 3044 3310 3045 3316
rect 3050 3311 3051 3316
rect 3074 3315 3075 3320
rect 3080 3315 3081 3320
rect 3103 3316 3104 3321
rect 3109 3319 3110 3321
rect 3129 3319 3136 3320
rect 3209 3319 3216 3320
rect 3109 3316 3130 3319
rect 3103 3315 3130 3316
rect 3074 3314 3081 3315
rect 3104 3314 3130 3315
rect 3135 3314 3136 3319
rect 3075 3311 3080 3314
rect 3050 3310 3080 3311
rect 3044 3305 3080 3310
rect 3104 3288 3109 3314
rect 3129 3313 3136 3314
rect 3186 3314 3210 3319
rect 3215 3314 3216 3319
rect 2935 3282 3109 3288
rect 2935 3259 2940 3282
rect 2972 3260 3012 3261
rect 2934 3258 2941 3259
rect 2934 3253 2935 3258
rect 2940 3253 2941 3258
rect 2972 3256 3006 3260
rect 2934 3252 2941 3253
rect 2971 3255 2978 3256
rect 2971 3250 2972 3255
rect 2977 3250 2978 3255
rect 3005 3255 3006 3256
rect 3011 3255 3012 3260
rect 3044 3260 3080 3265
rect 3186 3263 3191 3314
rect 3209 3313 3216 3314
rect 3005 3254 3012 3255
rect 3029 3255 3036 3256
rect 2971 3249 2978 3250
rect 2982 3251 2989 3252
rect 2982 3246 2983 3251
rect 2988 3246 2989 3251
rect 3029 3250 3030 3255
rect 3035 3250 3036 3255
rect 3044 3254 3045 3260
rect 3050 3259 3080 3260
rect 3050 3254 3051 3259
rect 3075 3256 3080 3259
rect 3185 3262 3192 3263
rect 3185 3257 3186 3262
rect 3191 3257 3192 3262
rect 3185 3256 3192 3257
rect 3044 3253 3051 3254
rect 3074 3255 3081 3256
rect 3074 3250 3075 3255
rect 3080 3250 3081 3255
rect 3103 3254 3110 3255
rect 3029 3249 3036 3250
rect 3058 3249 3065 3250
rect 3074 3249 3081 3250
rect 3087 3249 3093 3250
rect 3030 3246 3035 3249
rect 2982 3241 3035 3246
rect 3058 3244 3059 3249
rect 3064 3244 3065 3249
rect 3087 3244 3088 3249
rect 3092 3244 3093 3249
rect 3058 3243 3093 3244
rect 3059 3239 3093 3243
rect 3103 3249 3104 3254
rect 3109 3249 3110 3254
rect 3103 3248 3110 3249
rect 3129 3248 3136 3249
rect 3103 3243 3130 3248
rect 3135 3243 3136 3248
rect 3248 3244 3253 3353
rect 3298 3315 3305 3316
rect 3298 3310 3299 3315
rect 3304 3310 3305 3315
rect 3298 3309 3305 3310
rect 3205 3243 3253 3244
rect 3103 3222 3108 3243
rect 3129 3242 3136 3243
rect 2936 3216 3108 3222
rect 3174 3238 3253 3243
rect 3299 3247 3304 3309
rect 3299 3241 3366 3247
rect 2936 3196 2941 3216
rect 2935 3195 2942 3196
rect 2935 3190 2936 3195
rect 2941 3190 2942 3195
rect 2935 3189 2942 3190
rect 2982 3192 3035 3197
rect 3059 3195 3093 3199
rect 3174 3195 3179 3238
rect 2971 3188 2978 3189
rect 2971 3183 2972 3188
rect 2977 3183 2978 3188
rect 2982 3187 2983 3192
rect 2988 3187 2989 3192
rect 3030 3189 3035 3192
rect 3058 3194 3093 3195
rect 3058 3189 3059 3194
rect 3064 3189 3065 3194
rect 3087 3189 3088 3194
rect 3092 3189 3093 3194
rect 3173 3194 3180 3195
rect 2982 3186 2989 3187
rect 3029 3188 3036 3189
rect 3058 3188 3065 3189
rect 3074 3188 3081 3189
rect 3087 3188 3093 3189
rect 3103 3189 3110 3190
rect 2971 3182 2978 3183
rect 3005 3183 3012 3184
rect 3005 3182 3006 3183
rect 2972 3178 3006 3182
rect 3011 3178 3012 3183
rect 3029 3183 3030 3188
rect 3035 3183 3036 3188
rect 3029 3182 3036 3183
rect 3044 3184 3051 3185
rect 2972 3177 3012 3178
rect 3044 3178 3045 3184
rect 3050 3179 3051 3184
rect 3074 3183 3075 3188
rect 3080 3183 3081 3188
rect 3103 3184 3104 3189
rect 3109 3184 3110 3189
rect 3173 3189 3174 3194
rect 3179 3189 3180 3194
rect 3243 3192 3296 3197
rect 3320 3195 3354 3199
rect 3361 3195 3366 3241
rect 3173 3188 3180 3189
rect 3232 3188 3239 3189
rect 3103 3183 3110 3184
rect 3128 3183 3135 3184
rect 3074 3182 3081 3183
rect 3075 3179 3080 3182
rect 3050 3178 3080 3179
rect 3044 3173 3080 3178
rect 3105 3178 3129 3183
rect 3134 3178 3135 3183
rect 3232 3183 3233 3188
rect 3238 3183 3239 3188
rect 3243 3187 3244 3192
rect 3249 3187 3250 3192
rect 3291 3189 3296 3192
rect 3319 3194 3354 3195
rect 3319 3189 3320 3194
rect 3325 3189 3326 3194
rect 3348 3189 3349 3194
rect 3353 3189 3354 3194
rect 3243 3186 3250 3187
rect 3290 3188 3297 3189
rect 3319 3188 3326 3189
rect 3335 3188 3342 3189
rect 3348 3188 3354 3189
rect 3360 3194 3367 3195
rect 3360 3189 3361 3194
rect 3366 3189 3367 3194
rect 3360 3188 3367 3189
rect 3232 3182 3239 3183
rect 3266 3183 3273 3184
rect 3266 3182 3267 3183
rect 3105 3047 3110 3178
rect 3128 3177 3135 3178
rect 3233 3178 3267 3182
rect 3272 3178 3273 3183
rect 3290 3183 3291 3188
rect 3296 3183 3297 3188
rect 3290 3182 3297 3183
rect 3305 3184 3312 3185
rect 3233 3177 3273 3178
rect 3305 3178 3306 3184
rect 3311 3179 3312 3184
rect 3335 3183 3336 3188
rect 3341 3183 3342 3188
rect 3335 3182 3342 3183
rect 3336 3179 3341 3182
rect 3311 3178 3341 3179
rect 3305 3173 3341 3178
rect 3388 3150 3393 3677
rect 3235 3145 3393 3150
rect 3235 3083 3240 3145
rect 3234 3082 3240 3083
rect 3234 3078 3235 3082
rect 3239 3078 3240 3082
rect 3234 3077 3240 3078
rect 3105 3041 3416 3047
rect 3359 3000 3365 3001
rect 3359 2996 3360 3000
rect 3364 2996 3365 3000
rect 3359 2995 3365 2996
rect 2160 2804 2915 2810
rect 3360 2791 3365 2995
rect 1507 2786 3365 2791
rect 1507 2213 1512 2786
rect 1901 2751 1992 2752
rect 1901 2747 1987 2751
rect 1991 2747 1992 2751
rect 1902 2716 1907 2747
rect 1986 2746 1992 2747
rect 2931 2751 2937 2752
rect 2931 2747 2932 2751
rect 2936 2747 2937 2751
rect 2931 2746 2937 2747
rect 1763 2715 1907 2716
rect 1763 2711 1764 2715
rect 1768 2711 1907 2715
rect 2708 2716 2714 2717
rect 2931 2716 2936 2746
rect 1763 2710 1769 2711
rect 1989 2708 2469 2713
rect 2708 2712 2709 2716
rect 2713 2712 2936 2716
rect 3411 2713 3416 3041
rect 2708 2711 2936 2712
rect 3074 2708 3416 2713
rect 1989 2673 1994 2708
rect 2464 2703 3102 2708
rect 2442 2700 2448 2701
rect 2442 2696 2443 2700
rect 2447 2696 2448 2700
rect 2442 2695 2448 2696
rect 3387 2700 3393 2701
rect 3387 2696 3388 2700
rect 3392 2696 3393 2700
rect 3387 2695 3393 2696
rect 2027 2674 2067 2675
rect 1988 2672 1995 2673
rect 1988 2667 1989 2672
rect 1994 2667 1995 2672
rect 2027 2670 2061 2674
rect 1988 2666 1995 2667
rect 2026 2669 2033 2670
rect 2026 2664 2027 2669
rect 2032 2664 2033 2669
rect 2060 2669 2061 2670
rect 2066 2669 2067 2674
rect 2099 2674 2135 2679
rect 2060 2668 2067 2669
rect 2084 2669 2091 2670
rect 2026 2663 2033 2664
rect 2037 2665 2044 2666
rect 2037 2660 2038 2665
rect 2043 2660 2044 2665
rect 2084 2664 2085 2669
rect 2090 2664 2091 2669
rect 2099 2668 2100 2674
rect 2105 2673 2135 2674
rect 2105 2668 2106 2673
rect 2130 2670 2135 2673
rect 2099 2667 2106 2668
rect 2129 2669 2136 2670
rect 2129 2664 2130 2669
rect 2135 2664 2136 2669
rect 2158 2668 2165 2669
rect 2084 2663 2091 2664
rect 2113 2663 2120 2664
rect 2129 2663 2136 2664
rect 2142 2663 2148 2664
rect 2085 2660 2090 2663
rect 2037 2655 2090 2660
rect 2113 2658 2114 2663
rect 2119 2658 2120 2663
rect 2142 2658 2143 2663
rect 2147 2658 2148 2663
rect 2113 2657 2148 2658
rect 2114 2653 2148 2657
rect 2158 2663 2159 2668
rect 2164 2663 2165 2668
rect 2240 2668 2247 2669
rect 2240 2663 2241 2668
rect 2246 2663 2247 2668
rect 2325 2668 2332 2669
rect 2325 2663 2326 2668
rect 2331 2663 2332 2668
rect 2158 2662 2165 2663
rect 2184 2662 2191 2663
rect 2240 2662 2247 2663
rect 2265 2662 2272 2663
rect 2325 2662 2332 2663
rect 2158 2657 2185 2662
rect 2190 2657 2191 2662
rect 2241 2657 2266 2662
rect 2271 2657 2272 2662
rect 2158 2636 2163 2657
rect 2184 2656 2191 2657
rect 2265 2656 2272 2657
rect 2322 2657 2331 2662
rect 1991 2630 2163 2636
rect 1762 2612 1768 2613
rect 1762 2608 1763 2612
rect 1767 2608 1900 2612
rect 1991 2610 1996 2630
rect 1762 2607 1900 2608
rect 1506 2212 1512 2213
rect 1506 2208 1507 2212
rect 1511 2208 1512 2212
rect 1506 2207 1512 2208
rect 1895 1846 1900 2607
rect 1990 2609 1997 2610
rect 1990 2604 1991 2609
rect 1996 2604 1997 2609
rect 1990 2603 1997 2604
rect 2037 2606 2090 2611
rect 2114 2609 2148 2613
rect 2026 2602 2033 2603
rect 2026 2597 2027 2602
rect 2032 2597 2033 2602
rect 2037 2601 2038 2606
rect 2043 2601 2044 2606
rect 2085 2603 2090 2606
rect 2113 2608 2148 2609
rect 2113 2603 2114 2608
rect 2119 2603 2120 2608
rect 2142 2603 2143 2608
rect 2147 2603 2148 2608
rect 2037 2600 2044 2601
rect 2084 2602 2091 2603
rect 2113 2602 2120 2603
rect 2129 2602 2136 2603
rect 2142 2602 2148 2603
rect 2158 2603 2165 2604
rect 2184 2603 2191 2604
rect 2264 2603 2271 2604
rect 2026 2596 2033 2597
rect 2060 2597 2067 2598
rect 2060 2596 2061 2597
rect 2027 2592 2061 2596
rect 2066 2592 2067 2597
rect 2084 2597 2085 2602
rect 2090 2597 2091 2602
rect 2084 2596 2091 2597
rect 2099 2598 2106 2599
rect 2027 2591 2067 2592
rect 2099 2592 2100 2598
rect 2105 2593 2106 2598
rect 2129 2597 2130 2602
rect 2135 2597 2136 2602
rect 2158 2598 2159 2603
rect 2164 2598 2185 2603
rect 2190 2598 2191 2603
rect 2158 2597 2165 2598
rect 2184 2597 2191 2598
rect 2241 2598 2265 2603
rect 2270 2598 2271 2603
rect 2129 2596 2136 2597
rect 2130 2593 2135 2596
rect 2105 2592 2135 2593
rect 2099 2587 2135 2592
rect 2159 2570 2164 2597
rect 1990 2564 2164 2570
rect 1990 2541 1995 2564
rect 2027 2542 2067 2543
rect 1989 2540 1996 2541
rect 1989 2535 1990 2540
rect 1995 2535 1996 2540
rect 2027 2538 2061 2542
rect 1989 2534 1996 2535
rect 2026 2537 2033 2538
rect 2026 2532 2027 2537
rect 2032 2532 2033 2537
rect 2060 2537 2061 2538
rect 2066 2537 2067 2542
rect 2099 2542 2135 2547
rect 2241 2545 2246 2598
rect 2264 2597 2271 2598
rect 2322 2569 2327 2657
rect 2284 2564 2327 2569
rect 2060 2536 2067 2537
rect 2084 2537 2091 2538
rect 2026 2531 2033 2532
rect 2037 2533 2044 2534
rect 2037 2528 2038 2533
rect 2043 2528 2044 2533
rect 2084 2532 2085 2537
rect 2090 2532 2091 2537
rect 2099 2536 2100 2542
rect 2105 2541 2135 2542
rect 2105 2536 2106 2541
rect 2130 2538 2135 2541
rect 2240 2544 2247 2545
rect 2240 2539 2241 2544
rect 2246 2539 2247 2544
rect 2240 2538 2247 2539
rect 2099 2535 2106 2536
rect 2129 2537 2136 2538
rect 2129 2532 2130 2537
rect 2135 2532 2136 2537
rect 2158 2536 2165 2537
rect 2084 2531 2091 2532
rect 2113 2531 2120 2532
rect 2129 2531 2136 2532
rect 2142 2531 2148 2532
rect 2085 2528 2090 2531
rect 2037 2523 2090 2528
rect 2113 2526 2114 2531
rect 2119 2526 2120 2531
rect 2142 2526 2143 2531
rect 2147 2526 2148 2531
rect 2113 2525 2148 2526
rect 2114 2521 2148 2525
rect 2158 2531 2159 2536
rect 2164 2531 2165 2536
rect 2284 2531 2289 2564
rect 2347 2541 2354 2542
rect 2347 2536 2348 2541
rect 2353 2536 2354 2541
rect 2347 2535 2354 2536
rect 2158 2530 2165 2531
rect 2184 2530 2191 2531
rect 2158 2525 2185 2530
rect 2190 2525 2191 2530
rect 2284 2530 2296 2531
rect 2284 2525 2290 2530
rect 2295 2525 2296 2530
rect 2158 2504 2163 2525
rect 2184 2524 2191 2525
rect 2289 2524 2296 2525
rect 1991 2498 2163 2504
rect 1991 2478 1996 2498
rect 1990 2477 1997 2478
rect 1990 2472 1991 2477
rect 1996 2472 1997 2477
rect 1990 2471 1997 2472
rect 2037 2474 2090 2479
rect 2114 2477 2148 2481
rect 2026 2470 2033 2471
rect 2026 2465 2027 2470
rect 2032 2465 2033 2470
rect 2037 2469 2038 2474
rect 2043 2469 2044 2474
rect 2085 2471 2090 2474
rect 2113 2476 2148 2477
rect 2113 2471 2114 2476
rect 2119 2471 2120 2476
rect 2142 2471 2143 2476
rect 2147 2471 2148 2476
rect 2183 2472 2190 2473
rect 2289 2472 2296 2473
rect 2037 2468 2044 2469
rect 2084 2470 2091 2471
rect 2113 2470 2120 2471
rect 2129 2470 2136 2471
rect 2142 2470 2148 2471
rect 2158 2471 2184 2472
rect 2026 2464 2033 2465
rect 2060 2465 2067 2466
rect 2060 2464 2061 2465
rect 2027 2460 2061 2464
rect 2066 2460 2067 2465
rect 2084 2465 2085 2470
rect 2090 2465 2091 2470
rect 2084 2464 2091 2465
rect 2099 2466 2106 2467
rect 2027 2459 2067 2460
rect 2099 2460 2100 2466
rect 2105 2461 2106 2466
rect 2129 2465 2130 2470
rect 2135 2465 2136 2470
rect 2129 2464 2136 2465
rect 2158 2466 2159 2471
rect 2164 2467 2184 2471
rect 2189 2467 2190 2472
rect 2164 2466 2165 2467
rect 2183 2466 2190 2467
rect 2285 2467 2290 2472
rect 2295 2467 2296 2472
rect 2285 2466 2296 2467
rect 2158 2465 2165 2466
rect 2130 2461 2135 2464
rect 2105 2460 2135 2461
rect 2099 2455 2135 2460
rect 2158 2438 2163 2465
rect 1990 2432 2163 2438
rect 2285 2438 2290 2466
rect 2285 2433 2328 2438
rect 1990 2409 1995 2432
rect 2027 2410 2067 2411
rect 1989 2408 1996 2409
rect 1989 2403 1990 2408
rect 1995 2403 1996 2408
rect 2027 2406 2061 2410
rect 1989 2402 1996 2403
rect 2026 2405 2033 2406
rect 2026 2400 2027 2405
rect 2032 2400 2033 2405
rect 2060 2405 2061 2406
rect 2066 2405 2067 2410
rect 2099 2410 2135 2415
rect 2323 2414 2328 2433
rect 2060 2404 2067 2405
rect 2084 2405 2091 2406
rect 2026 2399 2033 2400
rect 2037 2401 2044 2402
rect 2037 2396 2038 2401
rect 2043 2396 2044 2401
rect 2084 2400 2085 2405
rect 2090 2400 2091 2405
rect 2099 2404 2100 2410
rect 2105 2409 2135 2410
rect 2105 2404 2106 2409
rect 2130 2406 2135 2409
rect 2322 2413 2329 2414
rect 2322 2408 2323 2413
rect 2328 2408 2329 2413
rect 2322 2407 2329 2408
rect 2348 2406 2353 2535
rect 2356 2406 2363 2407
rect 2099 2403 2106 2404
rect 2129 2405 2136 2406
rect 2129 2400 2130 2405
rect 2135 2400 2136 2405
rect 2158 2404 2165 2405
rect 2084 2399 2091 2400
rect 2113 2399 2120 2400
rect 2129 2399 2136 2400
rect 2142 2399 2148 2400
rect 2085 2396 2090 2399
rect 2037 2391 2090 2396
rect 2113 2394 2114 2399
rect 2119 2394 2120 2399
rect 2142 2394 2143 2399
rect 2147 2394 2148 2399
rect 2113 2393 2148 2394
rect 2114 2389 2148 2393
rect 2158 2399 2159 2404
rect 2164 2399 2165 2404
rect 2240 2404 2247 2405
rect 2240 2399 2241 2404
rect 2246 2399 2247 2404
rect 2336 2401 2357 2406
rect 2362 2401 2363 2406
rect 2336 2400 2348 2401
rect 2356 2400 2363 2401
rect 2158 2398 2165 2399
rect 2184 2398 2191 2399
rect 2240 2398 2247 2399
rect 2265 2398 2272 2399
rect 2158 2393 2185 2398
rect 2190 2393 2191 2398
rect 2241 2393 2266 2398
rect 2271 2393 2272 2398
rect 2158 2372 2163 2393
rect 2184 2392 2191 2393
rect 2265 2392 2272 2393
rect 2336 2392 2341 2400
rect 1991 2366 2163 2372
rect 2303 2371 2341 2392
rect 1991 2346 1996 2366
rect 1990 2345 1997 2346
rect 1990 2340 1991 2345
rect 1996 2340 1997 2345
rect 1990 2339 1997 2340
rect 2037 2342 2090 2347
rect 2114 2345 2148 2349
rect 2026 2338 2033 2339
rect 2026 2333 2027 2338
rect 2032 2333 2033 2338
rect 2037 2337 2038 2342
rect 2043 2337 2044 2342
rect 2085 2339 2090 2342
rect 2113 2344 2148 2345
rect 2113 2339 2114 2344
rect 2119 2339 2120 2344
rect 2142 2339 2143 2344
rect 2147 2339 2148 2344
rect 2037 2336 2044 2337
rect 2084 2338 2091 2339
rect 2113 2338 2120 2339
rect 2129 2338 2136 2339
rect 2142 2338 2148 2339
rect 2158 2339 2165 2340
rect 2026 2332 2033 2333
rect 2060 2333 2067 2334
rect 2060 2332 2061 2333
rect 2027 2328 2061 2332
rect 2066 2328 2067 2333
rect 2084 2333 2085 2338
rect 2090 2333 2091 2338
rect 2084 2332 2091 2333
rect 2099 2334 2106 2335
rect 2027 2327 2067 2328
rect 2099 2328 2100 2334
rect 2105 2329 2106 2334
rect 2129 2333 2130 2338
rect 2135 2333 2136 2338
rect 2158 2334 2159 2339
rect 2164 2337 2165 2339
rect 2184 2337 2191 2338
rect 2264 2337 2271 2338
rect 2164 2334 2185 2337
rect 2158 2333 2185 2334
rect 2129 2332 2136 2333
rect 2159 2332 2185 2333
rect 2190 2332 2191 2337
rect 2130 2329 2135 2332
rect 2105 2328 2135 2329
rect 2099 2323 2135 2328
rect 2159 2306 2164 2332
rect 2184 2331 2191 2332
rect 2241 2332 2265 2337
rect 2270 2332 2271 2337
rect 1990 2300 2164 2306
rect 1990 2277 1995 2300
rect 2027 2278 2067 2279
rect 1989 2276 1996 2277
rect 1989 2271 1990 2276
rect 1995 2271 1996 2276
rect 2027 2274 2061 2278
rect 1989 2270 1996 2271
rect 2026 2273 2033 2274
rect 2026 2268 2027 2273
rect 2032 2268 2033 2273
rect 2060 2273 2061 2274
rect 2066 2273 2067 2278
rect 2099 2278 2135 2283
rect 2241 2281 2246 2332
rect 2264 2331 2271 2332
rect 2060 2272 2067 2273
rect 2084 2273 2091 2274
rect 2026 2267 2033 2268
rect 2037 2269 2044 2270
rect 2037 2264 2038 2269
rect 2043 2264 2044 2269
rect 2084 2268 2085 2273
rect 2090 2268 2091 2273
rect 2099 2272 2100 2278
rect 2105 2277 2135 2278
rect 2105 2272 2106 2277
rect 2130 2274 2135 2277
rect 2240 2280 2247 2281
rect 2240 2275 2241 2280
rect 2246 2275 2247 2280
rect 2240 2274 2247 2275
rect 2099 2271 2106 2272
rect 2129 2273 2136 2274
rect 2129 2268 2130 2273
rect 2135 2268 2136 2273
rect 2158 2272 2165 2273
rect 2084 2267 2091 2268
rect 2113 2267 2120 2268
rect 2129 2267 2136 2268
rect 2142 2267 2148 2268
rect 2085 2264 2090 2267
rect 2037 2259 2090 2264
rect 2113 2262 2114 2267
rect 2119 2262 2120 2267
rect 2142 2262 2143 2267
rect 2147 2262 2148 2267
rect 2113 2261 2148 2262
rect 2114 2257 2148 2261
rect 2158 2267 2159 2272
rect 2164 2267 2165 2272
rect 2158 2266 2165 2267
rect 2184 2266 2191 2267
rect 2158 2261 2185 2266
rect 2190 2261 2191 2266
rect 2303 2262 2308 2371
rect 2353 2333 2360 2334
rect 2353 2328 2354 2333
rect 2359 2328 2360 2333
rect 2353 2327 2360 2328
rect 2260 2261 2308 2262
rect 2158 2240 2163 2261
rect 2184 2260 2191 2261
rect 1991 2234 2163 2240
rect 2229 2256 2308 2261
rect 2354 2265 2359 2327
rect 2354 2259 2421 2265
rect 1991 2214 1996 2234
rect 1990 2213 1997 2214
rect 1990 2208 1991 2213
rect 1996 2208 1997 2213
rect 1990 2207 1997 2208
rect 2037 2210 2090 2215
rect 2114 2213 2148 2217
rect 2229 2213 2234 2256
rect 2026 2206 2033 2207
rect 2026 2201 2027 2206
rect 2032 2201 2033 2206
rect 2037 2205 2038 2210
rect 2043 2205 2044 2210
rect 2085 2207 2090 2210
rect 2113 2212 2148 2213
rect 2113 2207 2114 2212
rect 2119 2207 2120 2212
rect 2142 2207 2143 2212
rect 2147 2207 2148 2212
rect 2228 2212 2235 2213
rect 2037 2204 2044 2205
rect 2084 2206 2091 2207
rect 2113 2206 2120 2207
rect 2129 2206 2136 2207
rect 2142 2206 2148 2207
rect 2158 2207 2165 2208
rect 2026 2200 2033 2201
rect 2060 2201 2067 2202
rect 2060 2200 2061 2201
rect 2027 2196 2061 2200
rect 2066 2196 2067 2201
rect 2084 2201 2085 2206
rect 2090 2201 2091 2206
rect 2084 2200 2091 2201
rect 2099 2202 2106 2203
rect 2027 2195 2067 2196
rect 2099 2196 2100 2202
rect 2105 2197 2106 2202
rect 2129 2201 2130 2206
rect 2135 2201 2136 2206
rect 2158 2202 2159 2207
rect 2164 2202 2165 2207
rect 2228 2207 2229 2212
rect 2234 2207 2235 2212
rect 2298 2210 2351 2215
rect 2375 2213 2409 2217
rect 2416 2213 2421 2259
rect 2228 2206 2235 2207
rect 2287 2206 2294 2207
rect 2158 2201 2165 2202
rect 2183 2201 2190 2202
rect 2129 2200 2136 2201
rect 2130 2197 2135 2200
rect 2105 2196 2135 2197
rect 2099 2191 2135 2196
rect 2160 2196 2184 2201
rect 2189 2196 2190 2201
rect 2287 2201 2288 2206
rect 2293 2201 2294 2206
rect 2298 2205 2299 2210
rect 2304 2205 2305 2210
rect 2346 2207 2351 2210
rect 2374 2212 2409 2213
rect 2374 2207 2375 2212
rect 2380 2207 2381 2212
rect 2403 2207 2404 2212
rect 2408 2207 2409 2212
rect 2298 2204 2305 2205
rect 2345 2206 2352 2207
rect 2374 2206 2381 2207
rect 2390 2206 2397 2207
rect 2403 2206 2409 2207
rect 2415 2212 2422 2213
rect 2415 2207 2416 2212
rect 2421 2207 2422 2212
rect 2415 2206 2422 2207
rect 2287 2200 2294 2201
rect 2321 2201 2328 2202
rect 2321 2200 2322 2201
rect 1895 1845 1901 1846
rect 1895 1841 1896 1845
rect 1900 1841 1901 1845
rect 1895 1840 1901 1841
rect 2160 1843 2165 2196
rect 2183 2195 2190 2196
rect 2288 2196 2322 2200
rect 2327 2196 2328 2201
rect 2345 2201 2346 2206
rect 2351 2201 2352 2206
rect 2345 2200 2352 2201
rect 2360 2202 2367 2203
rect 2288 2195 2328 2196
rect 2360 2196 2361 2202
rect 2366 2197 2367 2202
rect 2390 2201 2391 2206
rect 2396 2201 2397 2206
rect 2390 2200 2397 2201
rect 2391 2197 2396 2200
rect 2366 2196 2396 2197
rect 2360 2191 2396 2196
rect 2443 2168 2448 2695
rect 2972 2674 3012 2675
rect 2933 2672 2940 2673
rect 2910 2667 2934 2672
rect 2939 2667 2940 2672
rect 2972 2670 3006 2674
rect 2707 2612 2713 2613
rect 2707 2608 2708 2612
rect 2712 2608 2845 2612
rect 2707 2607 2845 2608
rect 2451 2212 2457 2213
rect 2451 2208 2452 2212
rect 2456 2208 2457 2212
rect 2451 2207 2457 2208
rect 2290 2163 2448 2168
rect 2290 2101 2295 2163
rect 2289 2100 2295 2101
rect 2289 2096 2290 2100
rect 2294 2096 2295 2100
rect 2289 2095 2295 2096
rect 2452 2038 2457 2207
rect 2415 2033 2457 2038
rect 2415 2019 2420 2033
rect 2414 2018 2420 2019
rect 2414 2014 2415 2018
rect 2419 2014 2420 2018
rect 2414 2013 2420 2014
rect 2840 1846 2845 2607
rect 2840 1845 2846 1846
rect 2160 1838 2205 1843
rect 2840 1841 2841 1845
rect 2845 1841 2846 1845
rect 2840 1840 2846 1841
rect 2910 1834 2915 2667
rect 2933 2666 2940 2667
rect 2971 2669 2978 2670
rect 2971 2664 2972 2669
rect 2977 2664 2978 2669
rect 3005 2669 3006 2670
rect 3011 2669 3012 2674
rect 3044 2674 3080 2679
rect 3005 2668 3012 2669
rect 3029 2669 3036 2670
rect 2971 2663 2978 2664
rect 2982 2665 2989 2666
rect 2982 2660 2983 2665
rect 2988 2660 2989 2665
rect 3029 2664 3030 2669
rect 3035 2664 3036 2669
rect 3044 2668 3045 2674
rect 3050 2673 3080 2674
rect 3050 2668 3051 2673
rect 3075 2670 3080 2673
rect 3044 2667 3051 2668
rect 3074 2669 3081 2670
rect 3074 2664 3075 2669
rect 3080 2664 3081 2669
rect 3103 2668 3110 2669
rect 3029 2663 3036 2664
rect 3058 2663 3065 2664
rect 3074 2663 3081 2664
rect 3087 2663 3093 2664
rect 3030 2660 3035 2663
rect 2982 2655 3035 2660
rect 3058 2658 3059 2663
rect 3064 2658 3065 2663
rect 3087 2658 3088 2663
rect 3092 2658 3093 2663
rect 3058 2657 3093 2658
rect 3059 2653 3093 2657
rect 3103 2663 3104 2668
rect 3109 2663 3110 2668
rect 3185 2668 3192 2669
rect 3185 2663 3186 2668
rect 3191 2663 3192 2668
rect 3270 2668 3277 2669
rect 3270 2663 3271 2668
rect 3276 2663 3277 2668
rect 3103 2662 3110 2663
rect 3129 2662 3136 2663
rect 3185 2662 3192 2663
rect 3210 2662 3217 2663
rect 3270 2662 3277 2663
rect 3103 2657 3130 2662
rect 3135 2657 3136 2662
rect 3186 2657 3211 2662
rect 3216 2657 3217 2662
rect 3103 2636 3108 2657
rect 3129 2656 3136 2657
rect 3210 2656 3217 2657
rect 3267 2657 3276 2662
rect 2936 2630 3108 2636
rect 2936 2610 2941 2630
rect 2935 2609 2942 2610
rect 2935 2604 2936 2609
rect 2941 2604 2942 2609
rect 2935 2603 2942 2604
rect 2982 2606 3035 2611
rect 3059 2609 3093 2613
rect 2971 2602 2978 2603
rect 2971 2597 2972 2602
rect 2977 2597 2978 2602
rect 2982 2601 2983 2606
rect 2988 2601 2989 2606
rect 3030 2603 3035 2606
rect 3058 2608 3093 2609
rect 3058 2603 3059 2608
rect 3064 2603 3065 2608
rect 3087 2603 3088 2608
rect 3092 2603 3093 2608
rect 2982 2600 2989 2601
rect 3029 2602 3036 2603
rect 3058 2602 3065 2603
rect 3074 2602 3081 2603
rect 3087 2602 3093 2603
rect 3103 2603 3110 2604
rect 3129 2603 3136 2604
rect 3209 2603 3216 2604
rect 2971 2596 2978 2597
rect 3005 2597 3012 2598
rect 3005 2596 3006 2597
rect 2972 2592 3006 2596
rect 3011 2592 3012 2597
rect 3029 2597 3030 2602
rect 3035 2597 3036 2602
rect 3029 2596 3036 2597
rect 3044 2598 3051 2599
rect 2972 2591 3012 2592
rect 3044 2592 3045 2598
rect 3050 2593 3051 2598
rect 3074 2597 3075 2602
rect 3080 2597 3081 2602
rect 3103 2598 3104 2603
rect 3109 2598 3130 2603
rect 3135 2598 3136 2603
rect 3103 2597 3110 2598
rect 3129 2597 3136 2598
rect 3186 2598 3210 2603
rect 3215 2598 3216 2603
rect 3074 2596 3081 2597
rect 3075 2593 3080 2596
rect 3050 2592 3080 2593
rect 3044 2587 3080 2592
rect 3104 2570 3109 2597
rect 2935 2564 3109 2570
rect 2935 2541 2940 2564
rect 2972 2542 3012 2543
rect 2934 2540 2941 2541
rect 2934 2535 2935 2540
rect 2940 2535 2941 2540
rect 2972 2538 3006 2542
rect 2934 2534 2941 2535
rect 2971 2537 2978 2538
rect 2971 2532 2972 2537
rect 2977 2532 2978 2537
rect 3005 2537 3006 2538
rect 3011 2537 3012 2542
rect 3044 2542 3080 2547
rect 3186 2545 3191 2598
rect 3209 2597 3216 2598
rect 3267 2569 3272 2657
rect 3229 2564 3272 2569
rect 3005 2536 3012 2537
rect 3029 2537 3036 2538
rect 2971 2531 2978 2532
rect 2982 2533 2989 2534
rect 2982 2528 2983 2533
rect 2988 2528 2989 2533
rect 3029 2532 3030 2537
rect 3035 2532 3036 2537
rect 3044 2536 3045 2542
rect 3050 2541 3080 2542
rect 3050 2536 3051 2541
rect 3075 2538 3080 2541
rect 3185 2544 3192 2545
rect 3185 2539 3186 2544
rect 3191 2539 3192 2544
rect 3185 2538 3192 2539
rect 3044 2535 3051 2536
rect 3074 2537 3081 2538
rect 3074 2532 3075 2537
rect 3080 2532 3081 2537
rect 3103 2536 3110 2537
rect 3029 2531 3036 2532
rect 3058 2531 3065 2532
rect 3074 2531 3081 2532
rect 3087 2531 3093 2532
rect 3030 2528 3035 2531
rect 2982 2523 3035 2528
rect 3058 2526 3059 2531
rect 3064 2526 3065 2531
rect 3087 2526 3088 2531
rect 3092 2526 3093 2531
rect 3058 2525 3093 2526
rect 3059 2521 3093 2525
rect 3103 2531 3104 2536
rect 3109 2531 3110 2536
rect 3229 2531 3234 2564
rect 3292 2541 3299 2542
rect 3292 2536 3293 2541
rect 3298 2536 3299 2541
rect 3292 2535 3299 2536
rect 3103 2530 3110 2531
rect 3129 2530 3136 2531
rect 3103 2525 3130 2530
rect 3135 2525 3136 2530
rect 3229 2530 3241 2531
rect 3229 2525 3235 2530
rect 3240 2525 3241 2530
rect 3103 2504 3108 2525
rect 3129 2524 3136 2525
rect 3234 2524 3241 2525
rect 2936 2498 3108 2504
rect 2936 2478 2941 2498
rect 2935 2477 2942 2478
rect 2935 2472 2936 2477
rect 2941 2472 2942 2477
rect 2935 2471 2942 2472
rect 2982 2474 3035 2479
rect 3059 2477 3093 2481
rect 2971 2470 2978 2471
rect 2971 2465 2972 2470
rect 2977 2465 2978 2470
rect 2982 2469 2983 2474
rect 2988 2469 2989 2474
rect 3030 2471 3035 2474
rect 3058 2476 3093 2477
rect 3058 2471 3059 2476
rect 3064 2471 3065 2476
rect 3087 2471 3088 2476
rect 3092 2471 3093 2476
rect 3128 2472 3135 2473
rect 3234 2472 3241 2473
rect 2982 2468 2989 2469
rect 3029 2470 3036 2471
rect 3058 2470 3065 2471
rect 3074 2470 3081 2471
rect 3087 2470 3093 2471
rect 3103 2471 3129 2472
rect 2971 2464 2978 2465
rect 3005 2465 3012 2466
rect 3005 2464 3006 2465
rect 2972 2460 3006 2464
rect 3011 2460 3012 2465
rect 3029 2465 3030 2470
rect 3035 2465 3036 2470
rect 3029 2464 3036 2465
rect 3044 2466 3051 2467
rect 2972 2459 3012 2460
rect 3044 2460 3045 2466
rect 3050 2461 3051 2466
rect 3074 2465 3075 2470
rect 3080 2465 3081 2470
rect 3074 2464 3081 2465
rect 3103 2466 3104 2471
rect 3109 2467 3129 2471
rect 3134 2467 3135 2472
rect 3109 2466 3110 2467
rect 3128 2466 3135 2467
rect 3230 2467 3235 2472
rect 3240 2467 3241 2472
rect 3230 2466 3241 2467
rect 3103 2465 3110 2466
rect 3075 2461 3080 2464
rect 3050 2460 3080 2461
rect 3044 2455 3080 2460
rect 3103 2438 3108 2465
rect 2935 2432 3108 2438
rect 3230 2438 3235 2466
rect 3230 2433 3273 2438
rect 2935 2409 2940 2432
rect 2972 2410 3012 2411
rect 2934 2408 2941 2409
rect 2934 2403 2935 2408
rect 2940 2403 2941 2408
rect 2972 2406 3006 2410
rect 2934 2402 2941 2403
rect 2971 2405 2978 2406
rect 2971 2400 2972 2405
rect 2977 2400 2978 2405
rect 3005 2405 3006 2406
rect 3011 2405 3012 2410
rect 3044 2410 3080 2415
rect 3268 2414 3273 2433
rect 3005 2404 3012 2405
rect 3029 2405 3036 2406
rect 2971 2399 2978 2400
rect 2982 2401 2989 2402
rect 2982 2396 2983 2401
rect 2988 2396 2989 2401
rect 3029 2400 3030 2405
rect 3035 2400 3036 2405
rect 3044 2404 3045 2410
rect 3050 2409 3080 2410
rect 3050 2404 3051 2409
rect 3075 2406 3080 2409
rect 3267 2413 3274 2414
rect 3267 2408 3268 2413
rect 3273 2408 3274 2413
rect 3267 2407 3274 2408
rect 3293 2406 3298 2535
rect 3301 2406 3308 2407
rect 3044 2403 3051 2404
rect 3074 2405 3081 2406
rect 3074 2400 3075 2405
rect 3080 2400 3081 2405
rect 3103 2404 3110 2405
rect 3029 2399 3036 2400
rect 3058 2399 3065 2400
rect 3074 2399 3081 2400
rect 3087 2399 3093 2400
rect 3030 2396 3035 2399
rect 2982 2391 3035 2396
rect 3058 2394 3059 2399
rect 3064 2394 3065 2399
rect 3087 2394 3088 2399
rect 3092 2394 3093 2399
rect 3058 2393 3093 2394
rect 3059 2389 3093 2393
rect 3103 2399 3104 2404
rect 3109 2399 3110 2404
rect 3185 2404 3192 2405
rect 3185 2399 3186 2404
rect 3191 2399 3192 2404
rect 3281 2401 3302 2406
rect 3307 2401 3308 2406
rect 3281 2400 3293 2401
rect 3301 2400 3308 2401
rect 3103 2398 3110 2399
rect 3129 2398 3136 2399
rect 3185 2398 3192 2399
rect 3210 2398 3217 2399
rect 3103 2393 3130 2398
rect 3135 2393 3136 2398
rect 3186 2393 3211 2398
rect 3216 2393 3217 2398
rect 3103 2372 3108 2393
rect 3129 2392 3136 2393
rect 3210 2392 3217 2393
rect 3281 2392 3286 2400
rect 2936 2366 3108 2372
rect 3248 2371 3286 2392
rect 2936 2346 2941 2366
rect 2935 2345 2942 2346
rect 2935 2340 2936 2345
rect 2941 2340 2942 2345
rect 2935 2339 2942 2340
rect 2982 2342 3035 2347
rect 3059 2345 3093 2349
rect 2971 2338 2978 2339
rect 2971 2333 2972 2338
rect 2977 2333 2978 2338
rect 2982 2337 2983 2342
rect 2988 2337 2989 2342
rect 3030 2339 3035 2342
rect 3058 2344 3093 2345
rect 3058 2339 3059 2344
rect 3064 2339 3065 2344
rect 3087 2339 3088 2344
rect 3092 2339 3093 2344
rect 2982 2336 2989 2337
rect 3029 2338 3036 2339
rect 3058 2338 3065 2339
rect 3074 2338 3081 2339
rect 3087 2338 3093 2339
rect 3103 2339 3110 2340
rect 2971 2332 2978 2333
rect 3005 2333 3012 2334
rect 3005 2332 3006 2333
rect 2972 2328 3006 2332
rect 3011 2328 3012 2333
rect 3029 2333 3030 2338
rect 3035 2333 3036 2338
rect 3029 2332 3036 2333
rect 3044 2334 3051 2335
rect 2972 2327 3012 2328
rect 3044 2328 3045 2334
rect 3050 2329 3051 2334
rect 3074 2333 3075 2338
rect 3080 2333 3081 2338
rect 3103 2334 3104 2339
rect 3109 2337 3110 2339
rect 3129 2337 3136 2338
rect 3209 2337 3216 2338
rect 3109 2334 3130 2337
rect 3103 2333 3130 2334
rect 3074 2332 3081 2333
rect 3104 2332 3130 2333
rect 3135 2332 3136 2337
rect 3075 2329 3080 2332
rect 3050 2328 3080 2329
rect 3044 2323 3080 2328
rect 3104 2306 3109 2332
rect 3129 2331 3136 2332
rect 3186 2332 3210 2337
rect 3215 2332 3216 2337
rect 2935 2300 3109 2306
rect 2935 2277 2940 2300
rect 2972 2278 3012 2279
rect 2934 2276 2941 2277
rect 2934 2271 2935 2276
rect 2940 2271 2941 2276
rect 2972 2274 3006 2278
rect 2934 2270 2941 2271
rect 2971 2273 2978 2274
rect 2971 2268 2972 2273
rect 2977 2268 2978 2273
rect 3005 2273 3006 2274
rect 3011 2273 3012 2278
rect 3044 2278 3080 2283
rect 3186 2281 3191 2332
rect 3209 2331 3216 2332
rect 3005 2272 3012 2273
rect 3029 2273 3036 2274
rect 2971 2267 2978 2268
rect 2982 2269 2989 2270
rect 2982 2264 2983 2269
rect 2988 2264 2989 2269
rect 3029 2268 3030 2273
rect 3035 2268 3036 2273
rect 3044 2272 3045 2278
rect 3050 2277 3080 2278
rect 3050 2272 3051 2277
rect 3075 2274 3080 2277
rect 3185 2280 3192 2281
rect 3185 2275 3186 2280
rect 3191 2275 3192 2280
rect 3185 2274 3192 2275
rect 3044 2271 3051 2272
rect 3074 2273 3081 2274
rect 3074 2268 3075 2273
rect 3080 2268 3081 2273
rect 3103 2272 3110 2273
rect 3029 2267 3036 2268
rect 3058 2267 3065 2268
rect 3074 2267 3081 2268
rect 3087 2267 3093 2268
rect 3030 2264 3035 2267
rect 2982 2259 3035 2264
rect 3058 2262 3059 2267
rect 3064 2262 3065 2267
rect 3087 2262 3088 2267
rect 3092 2262 3093 2267
rect 3058 2261 3093 2262
rect 3059 2257 3093 2261
rect 3103 2267 3104 2272
rect 3109 2267 3110 2272
rect 3103 2266 3110 2267
rect 3129 2266 3136 2267
rect 3103 2261 3130 2266
rect 3135 2261 3136 2266
rect 3248 2262 3253 2371
rect 3298 2333 3305 2334
rect 3298 2328 3299 2333
rect 3304 2328 3305 2333
rect 3298 2327 3305 2328
rect 3205 2261 3253 2262
rect 3103 2240 3108 2261
rect 3129 2260 3136 2261
rect 2936 2234 3108 2240
rect 3174 2256 3253 2261
rect 3299 2265 3304 2327
rect 3299 2259 3366 2265
rect 2936 2214 2941 2234
rect 2935 2213 2942 2214
rect 2935 2208 2936 2213
rect 2941 2208 2942 2213
rect 2935 2207 2942 2208
rect 2982 2210 3035 2215
rect 3059 2213 3093 2217
rect 3174 2213 3179 2256
rect 2971 2206 2978 2207
rect 2971 2201 2972 2206
rect 2977 2201 2978 2206
rect 2982 2205 2983 2210
rect 2988 2205 2989 2210
rect 3030 2207 3035 2210
rect 3058 2212 3093 2213
rect 3058 2207 3059 2212
rect 3064 2207 3065 2212
rect 3087 2207 3088 2212
rect 3092 2207 3093 2212
rect 3173 2212 3180 2213
rect 2982 2204 2989 2205
rect 3029 2206 3036 2207
rect 3058 2206 3065 2207
rect 3074 2206 3081 2207
rect 3087 2206 3093 2207
rect 3103 2207 3110 2208
rect 2971 2200 2978 2201
rect 3005 2201 3012 2202
rect 3005 2200 3006 2201
rect 2972 2196 3006 2200
rect 3011 2196 3012 2201
rect 3029 2201 3030 2206
rect 3035 2201 3036 2206
rect 3029 2200 3036 2201
rect 3044 2202 3051 2203
rect 2972 2195 3012 2196
rect 3044 2196 3045 2202
rect 3050 2197 3051 2202
rect 3074 2201 3075 2206
rect 3080 2201 3081 2206
rect 3103 2202 3104 2207
rect 3109 2202 3110 2207
rect 3173 2207 3174 2212
rect 3179 2207 3180 2212
rect 3243 2210 3296 2215
rect 3320 2213 3354 2217
rect 3361 2213 3366 2259
rect 3173 2206 3180 2207
rect 3232 2206 3239 2207
rect 3103 2201 3110 2202
rect 3128 2201 3135 2202
rect 3074 2200 3081 2201
rect 3075 2197 3080 2200
rect 3050 2196 3080 2197
rect 3105 2196 3129 2201
rect 3134 2196 3135 2201
rect 3232 2201 3233 2206
rect 3238 2201 3239 2206
rect 3243 2205 3244 2210
rect 3249 2205 3250 2210
rect 3291 2207 3296 2210
rect 3319 2212 3354 2213
rect 3319 2207 3320 2212
rect 3325 2207 3326 2212
rect 3348 2207 3349 2212
rect 3353 2207 3354 2212
rect 3243 2204 3250 2205
rect 3290 2206 3297 2207
rect 3319 2206 3326 2207
rect 3335 2206 3342 2207
rect 3348 2206 3354 2207
rect 3360 2212 3367 2213
rect 3360 2207 3361 2212
rect 3366 2207 3367 2212
rect 3360 2206 3367 2207
rect 3232 2200 3239 2201
rect 3266 2201 3273 2202
rect 3266 2200 3267 2201
rect 3044 2191 3080 2196
rect 3128 2195 3135 2196
rect 3233 2196 3267 2200
rect 3272 2196 3273 2201
rect 3290 2201 3291 2206
rect 3296 2201 3297 2206
rect 3290 2200 3297 2201
rect 3305 2202 3312 2203
rect 3233 2195 3273 2196
rect 3305 2196 3306 2202
rect 3311 2197 3312 2202
rect 3335 2201 3336 2206
rect 3341 2201 3342 2206
rect 3335 2200 3342 2201
rect 3336 2197 3341 2200
rect 3311 2196 3341 2197
rect 3305 2191 3341 2196
rect 3388 2168 3393 2695
rect 3235 2163 3393 2168
rect 3406 2212 3462 2217
rect 3235 2101 3240 2163
rect 3234 2100 3240 2101
rect 3234 2096 3235 2100
rect 3239 2096 3240 2100
rect 3234 2095 3240 2096
rect 3406 2038 3411 2212
rect 3360 2033 3411 2038
rect 3360 2019 3365 2033
rect 3359 2018 3365 2019
rect 3359 2014 3360 2018
rect 3364 2014 3365 2018
rect 3359 2013 3365 2014
rect 2160 1829 2915 1834
use BlankPad  t0
timestamp 1006127261
transform 1 0 960 0 1 4368
box -11 -51 298 632
use GNDPad  t1
timestamp 1509371954
transform 1 0 1258 0 1 4352
box 0 -35 309 648
use InPad  t2
timestamp 1509371954
transform 1 0 1599 0 1 4683
box -32 -366 277 317
use InPad  t3
timestamp 1509371954
transform 1 0 1908 0 1 4683
box -32 -366 277 317
use InPad  t4
timestamp 1509371954
transform 1 0 2217 0 1 4683
box -32 -366 277 317
use InPad  InPad_0
timestamp 1509371954
transform 1 0 2526 0 1 4683
box -32 -366 277 317
use InPad  InPad_1
timestamp 1509371954
transform 1 0 2835 0 1 4683
box -32 -366 277 317
use GNDPad  GNDPad_0
timestamp 1509371954
transform 1 0 3112 0 1 4352
box 0 -35 309 648
use VddPad  t8
timestamp 1509371954
transform 1 0 3421 0 1 4352
box 0 -35 309 648
use InPad  InPad_2
timestamp 1509371954
transform 1 0 3762 0 1 4683
box -32 -366 277 317
use Corner  crt
timestamp 1012241868
transform 0 1 4369 -1 0 4825
box -143 -333 774 618
use Corner  clt
timestamp 1012241868
transform 1 0 175 0 1 4369
box -143 -333 774 618
use BlankPad  l9
timestamp 1006127261
transform 0 -1 632 1 0 3740
box -11 -51 298 632
use BlankPad  l8
timestamp 1006127261
transform 0 -1 632 1 0 3431
box -11 -51 298 632
use BlankPad  l7
timestamp 1006127261
transform 0 -1 632 1 0 3122
box -11 -51 298 632
use BlankPad  l6
timestamp 1006127261
transform 0 -1 632 1 0 2813
box -11 -51 298 632
use BlankPad  l5
timestamp 1006127261
transform 0 -1 632 1 0 2504
box -11 -51 298 632
use BlankPad  l4
timestamp 1006127261
transform 0 -1 632 1 0 2195
box -11 -51 298 632
use BlankPad  l3
timestamp 1006127261
transform 0 -1 632 1 0 1886
box -11 -51 298 632
use BlankPad  l2
timestamp 1006127261
transform 0 -1 632 1 0 1577
box -11 -51 298 632
use BlankPad  l1
timestamp 1006127261
transform 0 -1 632 1 0 1268
box -11 -51 298 632
use BlankPad  r9
timestamp 1006127261
transform 0 1 4368 -1 0 4040
box -11 -51 298 632
use BlankPad  r8
timestamp 1006127261
transform 0 1 4368 -1 0 3731
box -11 -51 298 632
use BlankPad  r7
timestamp 1006127261
transform 0 1 4368 -1 0 3422
box -11 -51 298 632
use BlankPad  r6
timestamp 1006127261
transform 0 1 4368 -1 0 3113
box -11 -51 298 632
use BlankPad  r5
timestamp 1006127261
transform 0 1 4368 -1 0 2804
box -11 -51 298 632
use OutPad  OutPad_0
timestamp 1012172318
transform 0 1 4343 -1 0 2523
box 17 -26 326 657
use BlankPad  r3
timestamp 1006127261
transform 0 1 4368 -1 0 2186
box -11 -51 298 632
use BlankPad  r2
timestamp 1006127261
transform 0 1 4368 -1 0 1877
box -11 -51 298 632
use BlankPad  r1
timestamp 1006127261
transform 0 1 4368 -1 0 1568
box -11 -51 298 632
use BlankPad  r0
timestamp 1006127261
transform 0 1 4368 -1 0 1259
box -11 -51 298 632
use BlankPad  l0
timestamp 1006127261
transform 0 -1 632 1 0 959
box -11 -51 298 632
use Corner  clb
timestamp 1012241868
transform 0 -1 631 1 0 175
box -143 -333 774 618
use BlankPad  b0
timestamp 1006127261
transform -1 0 1260 0 -1 632
box -11 -51 298 632
use BlankPad  b1
timestamp 1006127261
transform -1 0 1569 0 -1 632
box -11 -51 298 632
use BlankPad  b2
timestamp 1006127261
transform -1 0 1878 0 -1 632
box -11 -51 298 632
use BlankPad  b3
timestamp 1006127261
transform -1 0 2187 0 -1 632
box -11 -51 298 632
use BlankPad  b4
timestamp 1006127261
transform -1 0 2496 0 -1 632
box -11 -51 298 632
use BlankPad  b5
timestamp 1006127261
transform -1 0 2805 0 -1 632
box -11 -51 298 632
use BlankPad  b6
timestamp 1006127261
transform -1 0 3114 0 -1 632
box -11 -51 298 632
use BlankPad  b7
timestamp 1006127261
transform -1 0 3423 0 -1 632
box -11 -51 298 632
use BlankPad  b8
timestamp 1006127261
transform -1 0 3732 0 -1 632
box -11 -51 298 632
use Corner  crb
timestamp 1012241868
transform -1 0 4825 0 -1 631
box -143 -333 774 618
use BlankPad  b9
timestamp 1006127261
transform -1 0 4041 0 -1 632
box -11 -51 298 632
<< labels >>
rlabel space 3809 4812 3953 4925 1 rst_b
rlabel metal1 3247 4840 3276 4906 1 GND!
rlabel metal1 2938 4844 2978 4893 1 mode
rlabel metal1 2629 4844 2669 4893 1 clk
rlabel metal1 2323 4847 2363 4896 1 data
rlabel metal1 2002 4848 2042 4897 1 program
rlabel space 4848 2311 4906 2362 1 out
rlabel metal1 3559 4267 3597 4306 1 Vdd!
rlabel metal1 2967 4285 2969 4288 1 Vdd!
<< end >>
