magic
tech scmos
timestamp 1607759597
<< ntransistor >>
rect 12 23 14 27
rect 28 23 30 27
rect 44 23 46 27
rect 67 23 69 27
rect 72 23 74 27
rect 98 23 100 27
rect 119 23 121 27
rect 139 23 141 27
rect 144 23 146 27
rect 162 23 164 27
rect 178 23 180 27
rect 194 23 196 27
rect 210 23 212 27
rect 233 23 235 27
rect 238 23 240 27
rect 264 23 266 27
rect 285 23 287 27
rect 305 23 307 27
rect 310 23 312 27
rect 328 23 330 27
rect 344 23 346 27
rect 360 23 362 27
rect 376 23 378 27
rect 399 23 401 27
rect 404 23 406 27
rect 430 23 432 27
rect 451 23 453 27
rect 471 23 473 27
rect 476 23 478 27
rect 494 23 496 27
rect 510 23 512 27
rect 526 23 528 27
rect 542 23 544 27
rect 565 23 567 27
rect 570 23 572 27
rect 596 23 598 27
rect 617 23 619 27
rect 637 23 639 27
rect 642 23 644 27
rect 660 23 662 27
<< ptransistor >>
rect 12 41 14 49
rect 28 41 30 49
rect 44 41 46 49
rect 67 41 69 49
rect 72 41 74 49
rect 98 41 100 49
rect 119 41 121 49
rect 139 41 141 49
rect 144 41 146 49
rect 162 41 164 49
rect 178 41 180 49
rect 194 41 196 49
rect 210 41 212 49
rect 233 41 235 49
rect 238 41 240 49
rect 264 41 266 49
rect 285 41 287 49
rect 305 41 307 49
rect 310 41 312 49
rect 328 41 330 49
rect 344 41 346 49
rect 360 41 362 49
rect 376 41 378 49
rect 399 41 401 49
rect 404 41 406 49
rect 430 41 432 49
rect 451 41 453 49
rect 471 41 473 49
rect 476 41 478 49
rect 494 41 496 49
rect 510 41 512 49
rect 526 41 528 49
rect 542 41 544 49
rect 565 41 567 49
rect 570 41 572 49
rect 596 41 598 49
rect 617 41 619 49
rect 637 41 639 49
rect 642 41 644 49
rect 660 41 662 49
<< ndiffusion >>
rect 11 23 12 27
rect 14 23 15 27
rect 27 23 28 27
rect 30 23 31 27
rect 43 23 44 27
rect 46 23 47 27
rect 62 23 67 27
rect 69 23 72 27
rect 74 23 75 27
rect 96 23 98 27
rect 100 23 101 27
rect 118 23 119 27
rect 121 23 122 27
rect 134 23 139 27
rect 141 23 144 27
rect 146 23 147 27
rect 161 23 162 27
rect 164 23 165 27
rect 177 23 178 27
rect 180 23 181 27
rect 193 23 194 27
rect 196 23 197 27
rect 209 23 210 27
rect 212 23 213 27
rect 228 23 233 27
rect 235 23 238 27
rect 240 23 241 27
rect 262 23 264 27
rect 266 23 267 27
rect 284 23 285 27
rect 287 23 288 27
rect 300 23 305 27
rect 307 23 310 27
rect 312 23 313 27
rect 327 23 328 27
rect 330 23 331 27
rect 343 23 344 27
rect 346 23 347 27
rect 359 23 360 27
rect 362 23 363 27
rect 375 23 376 27
rect 378 23 379 27
rect 394 23 399 27
rect 401 23 404 27
rect 406 23 407 27
rect 428 23 430 27
rect 432 23 433 27
rect 450 23 451 27
rect 453 23 454 27
rect 466 23 471 27
rect 473 23 476 27
rect 478 23 479 27
rect 493 23 494 27
rect 496 23 497 27
rect 509 23 510 27
rect 512 23 513 27
rect 525 23 526 27
rect 528 23 529 27
rect 541 23 542 27
rect 544 23 545 27
rect 560 23 565 27
rect 567 23 570 27
rect 572 23 573 27
rect 594 23 596 27
rect 598 23 599 27
rect 616 23 617 27
rect 619 23 620 27
rect 632 23 637 27
rect 639 23 642 27
rect 644 23 645 27
rect 659 23 660 27
rect 662 23 663 27
<< pdiffusion >>
rect 11 41 12 49
rect 14 41 15 49
rect 27 41 28 49
rect 30 41 31 49
rect 43 41 44 49
rect 46 41 47 49
rect 62 41 67 49
rect 69 41 72 49
rect 74 41 75 49
rect 96 41 98 49
rect 100 41 101 49
rect 118 41 119 49
rect 121 41 122 49
rect 134 41 139 49
rect 141 41 144 49
rect 146 41 147 49
rect 161 41 162 49
rect 164 41 165 49
rect 177 41 178 49
rect 180 41 181 49
rect 193 41 194 49
rect 196 41 197 49
rect 209 41 210 49
rect 212 41 213 49
rect 228 41 233 49
rect 235 41 238 49
rect 240 41 241 49
rect 262 41 264 49
rect 266 41 267 49
rect 284 41 285 49
rect 287 41 288 49
rect 300 41 305 49
rect 307 41 310 49
rect 312 41 313 49
rect 327 41 328 49
rect 330 41 331 49
rect 343 41 344 49
rect 346 41 347 49
rect 359 41 360 49
rect 362 41 363 49
rect 375 41 376 49
rect 378 41 379 49
rect 394 41 399 49
rect 401 41 404 49
rect 406 41 407 49
rect 428 41 430 49
rect 432 41 433 49
rect 450 41 451 49
rect 453 41 454 49
rect 466 41 471 49
rect 473 41 476 49
rect 478 41 479 49
rect 493 41 494 49
rect 496 41 497 49
rect 509 41 510 49
rect 512 41 513 49
rect 525 41 526 49
rect 528 41 529 49
rect 541 41 542 49
rect 544 41 545 49
rect 560 41 565 49
rect 567 41 570 49
rect 572 41 573 49
rect 594 41 596 49
rect 598 41 599 49
rect 616 41 617 49
rect 619 41 620 49
rect 632 41 637 49
rect 639 41 642 49
rect 644 41 645 49
rect 659 41 660 49
rect 662 41 663 49
<< ndcontact >>
rect 7 23 11 27
rect 15 23 19 27
rect 23 23 27 27
rect 31 23 35 27
rect 39 23 43 27
rect 47 23 51 27
rect 58 23 62 27
rect 75 23 79 27
rect 92 23 96 27
rect 101 23 105 27
rect 114 23 118 27
rect 122 23 126 27
rect 130 23 134 27
rect 147 23 151 27
rect 157 23 161 27
rect 165 23 169 27
rect 173 23 177 27
rect 181 23 185 27
rect 189 23 193 27
rect 197 23 201 27
rect 205 23 209 27
rect 213 23 217 27
rect 224 23 228 27
rect 241 23 245 27
rect 258 23 262 27
rect 267 23 271 27
rect 280 23 284 27
rect 288 23 292 27
rect 296 23 300 27
rect 313 23 317 27
rect 323 23 327 27
rect 331 23 335 27
rect 339 23 343 27
rect 347 23 351 27
rect 355 23 359 27
rect 363 23 367 27
rect 371 23 375 27
rect 379 23 383 27
rect 390 23 394 27
rect 407 23 411 27
rect 424 23 428 27
rect 433 23 437 27
rect 446 23 450 27
rect 454 23 458 27
rect 462 23 466 27
rect 479 23 483 27
rect 489 23 493 27
rect 497 23 501 27
rect 505 23 509 27
rect 513 23 517 27
rect 521 23 525 27
rect 529 23 533 27
rect 537 23 541 27
rect 545 23 549 27
rect 556 23 560 27
rect 573 23 577 27
rect 590 23 594 27
rect 599 23 603 27
rect 612 23 616 27
rect 620 23 624 27
rect 628 23 632 27
rect 645 23 649 27
rect 655 23 659 27
rect 663 23 667 27
<< pdcontact >>
rect 7 41 11 49
rect 15 41 19 49
rect 23 41 27 49
rect 31 41 35 49
rect 39 41 43 49
rect 47 41 51 49
rect 58 41 62 49
rect 75 41 79 49
rect 92 41 96 49
rect 101 41 105 49
rect 114 41 118 49
rect 122 41 126 49
rect 130 41 134 49
rect 147 41 151 49
rect 157 41 161 49
rect 165 41 169 49
rect 173 41 177 49
rect 181 41 185 49
rect 189 41 193 49
rect 197 41 201 49
rect 205 41 209 49
rect 213 41 217 49
rect 224 41 228 49
rect 241 41 245 49
rect 258 41 262 49
rect 267 41 271 49
rect 280 41 284 49
rect 288 41 292 49
rect 296 41 300 49
rect 313 41 317 49
rect 323 41 327 49
rect 331 41 335 49
rect 339 41 343 49
rect 347 41 351 49
rect 355 41 359 49
rect 363 41 367 49
rect 371 41 375 49
rect 379 41 383 49
rect 390 41 394 49
rect 407 41 411 49
rect 424 41 428 49
rect 433 41 437 49
rect 446 41 450 49
rect 454 41 458 49
rect 462 41 466 49
rect 479 41 483 49
rect 489 41 493 49
rect 497 41 501 49
rect 505 41 509 49
rect 513 41 517 49
rect 521 41 525 49
rect 529 41 533 49
rect 537 41 541 49
rect 545 41 549 49
rect 556 41 560 49
rect 573 41 577 49
rect 590 41 594 49
rect 599 41 603 49
rect 612 41 616 49
rect 620 41 624 49
rect 628 41 632 49
rect 645 41 649 49
rect 655 41 659 49
rect 663 41 667 49
<< psubstratepcontact >>
rect 0 7 4 11
rect 18 7 23 11
rect 48 7 52 11
rect 84 7 88 11
rect 123 7 127 11
rect 166 7 170 11
rect 184 7 189 11
rect 214 7 218 11
rect 250 7 254 11
rect 289 7 293 11
rect 332 7 336 11
rect 350 7 355 11
rect 380 7 384 11
rect 416 7 420 11
rect 455 7 459 11
rect 498 7 502 11
rect 516 7 521 11
rect 546 7 550 11
rect 582 7 586 11
rect 621 7 625 11
<< nsubstratencontact >>
rect 0 59 4 63
rect 18 59 23 63
rect 48 59 52 63
rect 84 59 88 63
rect 123 59 127 63
rect 166 59 170 63
rect 184 59 189 63
rect 214 59 218 63
rect 250 59 254 63
rect 289 59 293 63
rect 332 59 336 63
rect 350 59 355 63
rect 380 59 384 63
rect 416 59 420 63
rect 455 59 459 63
rect 498 59 502 63
rect 516 59 521 63
rect 546 59 550 63
rect 582 59 586 63
rect 621 59 625 63
<< polysilicon >>
rect 28 56 30 59
rect 72 56 74 59
rect 98 56 100 59
rect 144 56 146 59
rect 194 56 196 59
rect 238 56 240 59
rect 264 56 266 59
rect 310 56 312 59
rect 360 56 362 59
rect 404 56 406 59
rect 430 56 432 59
rect 476 56 478 59
rect 526 56 528 59
rect 570 56 572 59
rect 596 56 598 59
rect 642 56 644 59
rect 98 52 99 56
rect 264 52 265 56
rect 430 52 431 56
rect 596 52 597 56
rect 12 49 14 51
rect 28 49 30 52
rect 44 49 46 51
rect 67 49 69 51
rect 72 49 74 52
rect 98 49 100 52
rect 119 49 121 52
rect 139 49 141 51
rect 144 49 146 52
rect 162 49 164 51
rect 178 49 180 51
rect 194 49 196 52
rect 210 49 212 51
rect 233 49 235 51
rect 238 49 240 52
rect 264 49 266 52
rect 285 49 287 52
rect 305 49 307 51
rect 310 49 312 52
rect 328 49 330 51
rect 344 49 346 51
rect 360 49 362 52
rect 376 49 378 51
rect 399 49 401 51
rect 404 49 406 52
rect 430 49 432 52
rect 451 49 453 52
rect 471 49 473 51
rect 476 49 478 52
rect 494 49 496 51
rect 510 49 512 51
rect 526 49 528 52
rect 542 49 544 51
rect 565 49 567 51
rect 570 49 572 52
rect 596 49 598 52
rect 617 49 619 52
rect 637 49 639 51
rect 642 49 644 52
rect 660 49 662 51
rect 12 27 14 41
rect 28 39 30 41
rect 28 27 30 29
rect 44 27 46 41
rect 67 36 69 41
rect 72 39 74 41
rect 98 39 100 41
rect 63 32 69 36
rect 67 27 69 32
rect 72 27 74 29
rect 98 27 100 29
rect 119 27 121 41
rect 139 36 141 41
rect 144 39 146 41
rect 135 32 141 36
rect 139 27 141 32
rect 144 27 146 29
rect 162 27 164 41
rect 178 27 180 41
rect 194 39 196 41
rect 194 27 196 29
rect 210 27 212 41
rect 233 36 235 41
rect 238 39 240 41
rect 264 39 266 41
rect 229 32 235 36
rect 233 27 235 32
rect 238 27 240 29
rect 264 27 266 29
rect 285 27 287 41
rect 305 36 307 41
rect 310 39 312 41
rect 301 32 307 36
rect 305 27 307 32
rect 310 27 312 29
rect 328 27 330 41
rect 344 27 346 41
rect 360 39 362 41
rect 360 27 362 29
rect 376 27 378 41
rect 399 36 401 41
rect 404 39 406 41
rect 430 39 432 41
rect 395 32 401 36
rect 399 27 401 32
rect 404 27 406 29
rect 430 27 432 29
rect 451 27 453 41
rect 471 36 473 41
rect 476 39 478 41
rect 467 32 473 36
rect 471 27 473 32
rect 476 27 478 29
rect 494 27 496 41
rect 510 27 512 41
rect 526 39 528 41
rect 526 27 528 29
rect 542 27 544 41
rect 565 36 567 41
rect 570 39 572 41
rect 596 39 598 41
rect 561 32 567 36
rect 565 27 567 32
rect 570 27 572 29
rect 596 27 598 29
rect 617 27 619 41
rect 637 36 639 41
rect 642 39 644 41
rect 633 32 639 36
rect 637 27 639 32
rect 642 27 644 29
rect 660 27 662 41
rect 12 21 14 23
rect 28 19 30 23
rect 44 21 46 23
rect 67 21 69 23
rect 29 15 30 19
rect 72 18 74 23
rect 98 19 100 23
rect 119 21 121 23
rect 139 21 141 23
rect 28 12 30 15
rect 73 14 74 18
rect 99 15 100 19
rect 144 18 146 23
rect 162 21 164 23
rect 178 21 180 23
rect 194 19 196 23
rect 210 21 212 23
rect 233 21 235 23
rect 72 12 74 14
rect 98 11 100 15
rect 145 14 146 18
rect 195 15 196 19
rect 238 18 240 23
rect 264 19 266 23
rect 285 21 287 23
rect 305 21 307 23
rect 144 12 146 14
rect 194 12 196 15
rect 239 14 240 18
rect 265 15 266 19
rect 310 18 312 23
rect 328 21 330 23
rect 344 21 346 23
rect 360 19 362 23
rect 376 21 378 23
rect 399 21 401 23
rect 238 12 240 14
rect 264 11 266 15
rect 311 14 312 18
rect 361 15 362 19
rect 404 18 406 23
rect 430 19 432 23
rect 451 21 453 23
rect 471 21 473 23
rect 310 12 312 14
rect 360 12 362 15
rect 405 14 406 18
rect 431 15 432 19
rect 476 18 478 23
rect 494 21 496 23
rect 510 21 512 23
rect 526 19 528 23
rect 542 21 544 23
rect 565 21 567 23
rect 404 12 406 14
rect 430 11 432 15
rect 477 14 478 18
rect 527 15 528 19
rect 570 18 572 23
rect 596 19 598 23
rect 617 21 619 23
rect 637 21 639 23
rect 476 12 478 14
rect 526 12 528 15
rect 571 14 572 18
rect 597 15 598 19
rect 642 18 644 23
rect 660 21 662 23
rect 570 12 572 14
rect 596 11 598 15
rect 643 14 644 18
rect 642 12 644 14
<< polycontact >>
rect 28 52 32 56
rect 72 52 76 56
rect 99 52 103 56
rect 144 52 148 56
rect 194 52 198 56
rect 238 52 242 56
rect 265 52 269 56
rect 310 52 314 56
rect 360 52 364 56
rect 404 52 408 56
rect 431 52 435 56
rect 476 52 480 56
rect 526 52 530 56
rect 570 52 574 56
rect 597 52 601 56
rect 642 52 646 56
rect 8 32 12 36
rect 40 33 44 37
rect 59 32 63 36
rect 115 33 119 37
rect 131 32 135 36
rect 158 32 162 36
rect 174 32 178 36
rect 206 33 210 37
rect 225 32 229 36
rect 281 33 285 37
rect 297 32 301 36
rect 324 32 328 36
rect 340 32 344 36
rect 372 33 376 37
rect 391 32 395 36
rect 447 33 451 37
rect 463 32 467 36
rect 490 32 494 36
rect 506 32 510 36
rect 538 33 542 37
rect 557 32 561 36
rect 613 33 617 37
rect 629 32 633 36
rect 656 32 660 36
rect 25 15 29 19
rect 69 14 73 18
rect 94 15 99 19
rect 141 14 145 18
rect 191 15 195 19
rect 235 14 239 18
rect 260 15 265 19
rect 307 14 311 18
rect 357 15 361 19
rect 401 14 405 18
rect 426 15 431 19
rect 473 14 477 18
rect 523 15 527 19
rect 567 14 571 18
rect 592 15 597 19
rect 639 14 643 18
<< metal1 >>
rect 0 66 32 70
rect 36 66 61 70
rect 65 66 86 70
rect 90 66 150 70
rect 154 66 198 70
rect 202 66 227 70
rect 231 66 252 70
rect 256 66 316 70
rect 320 66 364 70
rect 368 66 393 70
rect 397 66 418 70
rect 422 66 482 70
rect 486 66 530 70
rect 534 66 559 70
rect 563 66 584 70
rect 588 66 648 70
rect 652 66 667 70
rect 4 59 18 63
rect 23 59 48 63
rect 52 59 84 63
rect 88 59 123 63
rect 127 59 166 63
rect 170 59 184 63
rect 189 59 214 63
rect 218 59 250 63
rect 254 59 289 63
rect 293 59 332 63
rect 336 59 350 63
rect 355 59 380 63
rect 384 59 416 63
rect 420 59 455 63
rect 459 59 498 63
rect 502 59 516 63
rect 521 59 546 63
rect 550 59 582 63
rect 586 59 621 63
rect 625 59 667 63
rect 7 49 10 59
rect 39 49 42 59
rect 58 49 61 59
rect 76 52 79 56
rect 103 52 104 56
rect 114 49 117 59
rect 130 49 133 59
rect 148 52 150 56
rect 157 49 160 59
rect 173 49 176 59
rect 205 49 208 59
rect 224 49 227 59
rect 242 52 245 56
rect 269 52 270 56
rect 280 49 283 59
rect 296 49 299 59
rect 314 52 316 56
rect 323 49 326 59
rect 339 49 342 59
rect 371 49 374 59
rect 390 49 393 59
rect 408 52 411 56
rect 435 52 436 56
rect 446 49 449 59
rect 462 49 465 59
rect 480 52 482 56
rect 489 49 492 59
rect 505 49 508 59
rect 537 49 540 59
rect 556 49 559 59
rect 574 52 577 56
rect 601 52 602 56
rect 612 49 615 59
rect 628 49 631 59
rect 646 52 648 56
rect 655 49 658 59
rect 3 32 8 35
rect 16 35 19 41
rect 23 35 26 41
rect 16 32 26 35
rect 16 27 19 32
rect 23 27 26 32
rect 32 37 35 41
rect 32 33 34 37
rect 38 33 40 37
rect 48 36 51 41
rect 76 38 79 41
rect 48 34 59 36
rect 32 27 35 33
rect 48 32 54 34
rect 48 27 51 32
rect 58 32 59 34
rect 77 34 79 38
rect 76 27 79 34
rect 92 37 95 41
rect 102 37 105 41
rect 102 33 111 37
rect 123 36 126 41
rect 148 37 151 41
rect 92 27 95 33
rect 102 27 105 33
rect 123 32 124 36
rect 128 32 131 35
rect 150 33 151 37
rect 123 27 126 32
rect 148 27 151 33
rect 166 35 169 41
rect 166 32 174 35
rect 182 35 185 41
rect 189 35 192 41
rect 182 32 192 35
rect 166 27 169 32
rect 182 27 185 32
rect 189 27 192 32
rect 198 37 201 41
rect 198 33 200 37
rect 204 33 206 37
rect 214 36 217 41
rect 242 38 245 41
rect 214 34 225 36
rect 198 27 201 33
rect 214 32 220 34
rect 214 27 217 32
rect 224 32 225 34
rect 243 34 245 38
rect 242 27 245 34
rect 258 37 261 41
rect 268 37 271 41
rect 268 33 277 37
rect 289 36 292 41
rect 314 37 317 41
rect 258 27 261 33
rect 268 27 271 33
rect 289 32 290 36
rect 294 32 297 35
rect 316 33 317 37
rect 289 27 292 32
rect 314 27 317 33
rect 332 35 335 41
rect 332 32 340 35
rect 348 35 351 41
rect 355 35 358 41
rect 348 32 358 35
rect 332 27 335 32
rect 348 27 351 32
rect 355 27 358 32
rect 364 37 367 41
rect 364 33 366 37
rect 370 33 372 37
rect 380 36 383 41
rect 408 38 411 41
rect 380 34 391 36
rect 364 27 367 33
rect 380 32 386 34
rect 380 27 383 32
rect 390 32 391 34
rect 409 34 411 38
rect 408 27 411 34
rect 424 37 427 41
rect 434 37 437 41
rect 434 33 443 37
rect 455 36 458 41
rect 480 37 483 41
rect 424 27 427 33
rect 434 27 437 33
rect 455 32 456 36
rect 460 32 463 35
rect 482 33 483 37
rect 455 27 458 32
rect 480 27 483 33
rect 498 35 501 41
rect 498 32 506 35
rect 514 35 517 41
rect 521 35 524 41
rect 514 32 524 35
rect 498 27 501 32
rect 514 27 517 32
rect 521 27 524 32
rect 530 37 533 41
rect 530 33 532 37
rect 536 33 538 37
rect 546 36 549 41
rect 574 38 577 41
rect 546 34 557 36
rect 530 27 533 33
rect 546 32 552 34
rect 546 27 549 32
rect 556 32 557 34
rect 575 34 577 38
rect 574 27 577 34
rect 590 37 593 41
rect 600 37 603 41
rect 600 33 609 37
rect 621 36 624 41
rect 646 37 649 41
rect 590 27 593 33
rect 600 27 603 33
rect 621 32 622 36
rect 626 32 629 35
rect 648 33 649 37
rect 621 27 624 32
rect 646 27 649 33
rect 664 27 667 41
rect 7 11 10 23
rect 39 11 42 23
rect 58 11 61 23
rect 68 14 69 18
rect 93 15 94 19
rect 114 11 117 23
rect 130 11 133 23
rect 140 14 141 18
rect 157 11 160 23
rect 173 11 176 23
rect 205 11 208 23
rect 224 11 227 23
rect 234 14 235 18
rect 259 15 260 19
rect 280 11 283 23
rect 296 11 299 23
rect 306 14 307 18
rect 323 11 326 23
rect 339 11 342 23
rect 371 11 374 23
rect 390 11 393 23
rect 400 14 401 18
rect 425 15 426 19
rect 446 11 449 23
rect 462 11 465 23
rect 472 14 473 18
rect 489 11 492 23
rect 505 11 508 23
rect 537 11 540 23
rect 556 11 559 23
rect 566 14 567 18
rect 591 15 592 19
rect 612 11 615 23
rect 628 11 631 23
rect 638 14 639 18
rect 655 11 658 23
rect 4 7 18 11
rect 23 7 48 11
rect 52 7 84 11
rect 88 7 123 11
rect 127 7 166 11
rect 170 7 184 11
rect 189 7 214 11
rect 218 7 250 11
rect 254 7 289 11
rect 293 7 332 11
rect 336 7 350 11
rect 355 7 380 11
rect 384 7 416 11
rect 420 7 455 11
rect 459 7 498 11
rect 502 7 516 11
rect 521 7 546 11
rect 550 7 582 11
rect 586 7 621 11
rect 625 7 667 11
rect 0 0 21 4
rect 25 0 80 4
rect 84 0 105 4
rect 109 0 136 4
rect 140 0 187 4
rect 191 0 246 4
rect 250 0 271 4
rect 275 0 302 4
rect 306 0 353 4
rect 357 0 412 4
rect 416 0 437 4
rect 441 0 468 4
rect 472 0 519 4
rect 523 0 578 4
rect 582 0 603 4
rect 607 0 634 4
rect 638 0 667 4
<< m2contact >>
rect 32 66 36 70
rect 61 66 65 70
rect 86 66 90 70
rect 150 66 154 70
rect 198 66 202 70
rect 227 66 231 70
rect 252 66 256 70
rect 316 66 320 70
rect 364 66 368 70
rect 393 66 397 70
rect 418 66 422 70
rect 482 66 486 70
rect 530 66 534 70
rect 559 66 563 70
rect 584 66 588 70
rect 648 66 652 70
rect 32 52 36 56
rect 79 52 83 56
rect 104 52 108 56
rect 150 52 154 56
rect 198 52 202 56
rect 245 52 249 56
rect 270 52 274 56
rect 316 52 320 56
rect 364 52 368 56
rect 411 52 415 56
rect 436 52 440 56
rect 482 52 486 56
rect 530 52 534 56
rect 577 52 581 56
rect 602 52 606 56
rect 648 52 652 56
rect 34 33 38 37
rect 54 30 58 34
rect 73 34 77 38
rect 92 33 96 37
rect 111 33 115 37
rect 124 32 128 36
rect 146 33 150 37
rect 154 32 158 36
rect 200 33 204 37
rect 220 30 224 34
rect 239 34 243 38
rect 258 33 262 37
rect 277 33 281 37
rect 290 32 294 36
rect 312 33 316 37
rect 320 32 324 36
rect 366 33 370 37
rect 386 30 390 34
rect 405 34 409 38
rect 424 33 428 37
rect 443 33 447 37
rect 456 32 460 36
rect 478 33 482 37
rect 486 32 490 36
rect 532 33 536 37
rect 552 30 556 34
rect 571 34 575 38
rect 590 33 594 37
rect 609 33 613 37
rect 622 32 626 36
rect 644 33 648 37
rect 652 32 656 36
rect 21 15 25 19
rect 64 14 68 18
rect 86 15 93 19
rect 136 14 140 18
rect 187 15 191 19
rect 230 14 234 18
rect 252 15 259 19
rect 302 14 306 18
rect 353 15 357 19
rect 396 14 400 18
rect 418 15 425 19
rect 468 14 472 18
rect 519 15 523 19
rect 562 14 566 18
rect 584 15 591 19
rect 634 14 638 18
rect 21 0 25 4
rect 80 0 84 4
rect 105 0 109 4
rect 136 0 140 4
rect 187 0 191 4
rect 246 0 250 4
rect 271 0 275 4
rect 302 0 306 4
rect 353 0 357 4
rect 412 0 416 4
rect 437 0 441 4
rect 468 0 472 4
rect 519 0 523 4
rect 578 0 582 4
rect 603 0 607 4
rect 634 0 638 4
<< metal2 >>
rect 33 56 36 66
rect 21 4 24 15
rect 61 14 64 66
rect 80 4 83 52
rect 86 19 89 66
rect 151 56 154 66
rect 199 56 202 66
rect 105 4 108 52
rect 136 4 140 14
rect 187 4 190 15
rect 227 14 230 66
rect 246 4 249 52
rect 252 19 255 66
rect 317 56 320 66
rect 365 56 368 66
rect 271 4 274 52
rect 302 4 306 14
rect 353 4 356 15
rect 393 14 396 66
rect 412 4 415 52
rect 418 19 421 66
rect 483 56 486 66
rect 531 56 534 66
rect 437 4 440 52
rect 468 4 472 14
rect 519 4 522 15
rect 559 14 562 66
rect 578 4 581 52
rect 584 19 587 66
rect 649 56 652 66
rect 603 4 606 52
rect 634 4 638 14
<< m3contact >>
rect 38 33 43 38
rect 53 25 58 30
rect 68 33 73 38
rect 96 33 101 38
rect 111 37 116 43
rect 141 33 146 38
rect 204 33 209 38
rect 125 27 130 32
rect 154 27 158 32
rect 219 25 224 30
rect 234 33 239 38
rect 262 33 267 38
rect 277 37 282 43
rect 307 33 312 38
rect 370 33 375 38
rect 291 27 296 32
rect 320 27 324 32
rect 385 25 390 30
rect 400 33 405 38
rect 428 33 433 38
rect 443 37 448 43
rect 473 33 478 38
rect 536 33 541 38
rect 457 27 462 32
rect 486 27 490 32
rect 551 25 556 30
rect 566 33 571 38
rect 594 33 599 38
rect 609 37 614 43
rect 639 33 644 38
rect 623 27 628 32
rect 652 27 656 32
<< metal3 >>
rect 38 39 73 44
rect 110 43 146 48
rect 37 38 44 39
rect 37 33 38 38
rect 43 33 44 38
rect 37 32 44 33
rect 67 38 74 39
rect 67 33 68 38
rect 73 33 74 38
rect 67 32 74 33
rect 95 38 102 39
rect 95 33 96 38
rect 101 33 102 38
rect 110 37 111 43
rect 116 42 146 43
rect 116 37 117 42
rect 141 39 146 42
rect 204 39 239 44
rect 276 43 312 48
rect 110 36 117 37
rect 140 38 147 39
rect 140 33 141 38
rect 146 33 147 38
rect 203 38 210 39
rect 203 33 204 38
rect 209 33 210 38
rect 95 32 102 33
rect 124 32 131 33
rect 140 32 147 33
rect 153 32 159 33
rect 203 32 210 33
rect 233 38 240 39
rect 233 33 234 38
rect 239 33 240 38
rect 233 32 240 33
rect 261 38 268 39
rect 261 33 262 38
rect 267 33 268 38
rect 276 37 277 43
rect 282 42 312 43
rect 282 37 283 42
rect 307 39 312 42
rect 370 39 405 44
rect 442 43 478 48
rect 276 36 283 37
rect 306 38 313 39
rect 306 33 307 38
rect 312 33 313 38
rect 369 38 376 39
rect 369 33 370 38
rect 375 33 376 38
rect 261 32 268 33
rect 290 32 297 33
rect 306 32 313 33
rect 319 32 325 33
rect 369 32 376 33
rect 399 38 406 39
rect 399 33 400 38
rect 405 33 406 38
rect 399 32 406 33
rect 427 38 434 39
rect 427 33 428 38
rect 433 33 434 38
rect 442 37 443 43
rect 448 42 478 43
rect 448 37 449 42
rect 473 39 478 42
rect 536 39 571 44
rect 608 43 644 48
rect 442 36 449 37
rect 472 38 479 39
rect 472 33 473 38
rect 478 33 479 38
rect 535 38 542 39
rect 535 33 536 38
rect 541 33 542 38
rect 427 32 434 33
rect 456 32 463 33
rect 472 32 479 33
rect 485 32 491 33
rect 535 32 542 33
rect 565 38 572 39
rect 565 33 566 38
rect 571 33 572 38
rect 565 32 572 33
rect 593 38 600 39
rect 593 33 594 38
rect 599 33 600 38
rect 608 37 609 43
rect 614 42 644 43
rect 614 37 615 42
rect 639 39 644 42
rect 608 36 615 37
rect 638 38 645 39
rect 638 33 639 38
rect 644 33 645 38
rect 593 32 600 33
rect 622 32 629 33
rect 638 32 645 33
rect 651 32 657 33
rect 52 30 59 31
rect 52 25 53 30
rect 58 29 59 30
rect 96 29 101 32
rect 58 25 101 29
rect 124 27 125 32
rect 130 27 131 32
rect 153 27 154 32
rect 158 27 159 32
rect 124 26 159 27
rect 52 24 101 25
rect 125 22 159 26
rect 218 30 225 31
rect 218 25 219 30
rect 224 29 225 30
rect 262 29 267 32
rect 224 25 267 29
rect 290 27 291 32
rect 296 27 297 32
rect 319 27 320 32
rect 324 27 325 32
rect 290 26 325 27
rect 218 24 267 25
rect 291 22 325 26
rect 384 30 391 31
rect 384 25 385 30
rect 390 29 391 30
rect 428 29 433 32
rect 390 25 433 29
rect 456 27 457 32
rect 462 27 463 32
rect 485 27 486 32
rect 490 27 491 32
rect 456 26 491 27
rect 384 24 433 25
rect 457 22 491 26
rect 550 30 557 31
rect 550 25 551 30
rect 556 29 557 30
rect 594 29 599 32
rect 556 25 599 29
rect 622 27 623 32
rect 628 27 629 32
rect 651 27 652 32
rect 656 27 657 32
rect 622 26 657 27
rect 550 24 599 25
rect 623 22 657 26
<< labels >>
rlabel metal1 3 32 7 35 1 D
rlabel metal1 8 7 11 11 1 GND!
rlabel metal1 7 59 10 63 1 Vdd!
rlabel metal1 0 66 3 70 4 clk
rlabel metal1 0 0 3 4 2 ~clk
rlabel metal1 166 0 169 4 2 ~clk
rlabel metal1 166 66 169 70 4 clk
rlabel metal1 173 59 176 63 1 Vdd!
rlabel metal1 174 7 177 11 1 GND!
rlabel metal1 169 32 173 35 1 q0
rlabel metal1 506 7 509 11 1 GND!
rlabel metal1 505 59 508 63 1 Vdd!
rlabel metal1 498 66 501 70 4 clk
rlabel metal1 498 0 501 4 2 ~clk
rlabel metal1 332 0 335 4 2 ~clk
rlabel metal1 332 66 335 70 4 clk
rlabel metal1 339 59 342 63 1 Vdd!
rlabel metal1 340 7 343 11 1 GND!
rlabel metal1 335 32 339 35 1 q1
rlabel metal1 501 32 505 35 1 q2
rlabel metal1 664 33 667 36 7 q3
<< end >>
