magic
tech scmos
timestamp 1608104755
<< ntransistor >>
rect 101 191 103 195
rect 106 191 108 195
rect 122 191 124 195
rect 138 191 140 195
rect 143 191 145 195
rect 164 191 166 195
rect 180 191 182 195
rect 196 191 198 195
rect 201 191 203 195
rect 217 191 219 195
rect 233 191 235 195
rect 238 191 240 195
rect 254 191 256 195
rect 270 191 272 195
rect 275 191 277 195
rect 296 191 298 195
rect 312 191 314 195
rect 328 191 330 195
rect 333 191 335 195
rect 349 191 351 195
rect 365 191 367 195
rect 370 191 372 195
rect 386 191 388 195
rect 402 191 404 195
rect 407 191 409 195
rect 428 191 430 195
rect 444 191 446 195
rect 460 191 462 195
rect 465 191 467 195
rect 481 191 483 195
<< ptransistor >>
rect 101 214 103 222
rect 106 214 108 222
rect 122 214 124 222
rect 138 214 140 222
rect 143 214 145 222
rect 164 214 166 222
rect 180 214 182 222
rect 196 214 198 222
rect 201 214 203 222
rect 217 214 219 222
rect 233 214 235 222
rect 238 214 240 222
rect 254 214 256 222
rect 270 214 272 222
rect 275 214 277 222
rect 296 214 298 222
rect 312 214 314 222
rect 328 214 330 222
rect 333 214 335 222
rect 349 214 351 222
rect 365 214 367 222
rect 370 214 372 222
rect 386 214 388 222
rect 402 214 404 222
rect 407 214 409 222
rect 428 214 430 222
rect 444 214 446 222
rect 460 214 462 222
rect 465 214 467 222
rect 481 214 483 222
<< ndiffusion >>
rect 100 191 101 195
rect 103 191 106 195
rect 108 191 109 195
rect 121 191 122 195
rect 124 191 125 195
rect 137 191 138 195
rect 140 191 143 195
rect 145 191 146 195
rect 163 191 164 195
rect 166 191 167 195
rect 179 191 180 195
rect 182 191 183 195
rect 195 191 196 195
rect 198 191 201 195
rect 203 191 204 195
rect 216 191 217 195
rect 219 191 220 195
rect 232 191 233 195
rect 235 191 238 195
rect 240 191 241 195
rect 253 191 254 195
rect 256 191 257 195
rect 269 191 270 195
rect 272 191 275 195
rect 277 191 278 195
rect 295 191 296 195
rect 298 191 299 195
rect 311 191 312 195
rect 314 191 315 195
rect 327 191 328 195
rect 330 191 333 195
rect 335 191 336 195
rect 348 191 349 195
rect 351 191 352 195
rect 364 191 365 195
rect 367 191 370 195
rect 372 191 373 195
rect 385 191 386 195
rect 388 191 389 195
rect 401 191 402 195
rect 404 191 407 195
rect 409 191 410 195
rect 427 191 428 195
rect 430 191 431 195
rect 443 191 444 195
rect 446 191 447 195
rect 459 191 460 195
rect 462 191 465 195
rect 467 191 468 195
rect 480 191 481 195
rect 483 191 484 195
<< pdiffusion >>
rect 100 214 101 222
rect 103 214 106 222
rect 108 214 109 222
rect 121 214 122 222
rect 124 218 125 222
rect 124 214 129 218
rect 137 214 138 222
rect 140 214 143 222
rect 145 214 146 222
rect 163 214 164 222
rect 166 214 167 222
rect 179 214 180 222
rect 182 218 183 222
rect 182 214 187 218
rect 195 214 196 222
rect 198 214 201 222
rect 203 214 204 222
rect 216 214 217 222
rect 219 214 220 222
rect 232 214 233 222
rect 235 214 238 222
rect 240 214 241 222
rect 253 214 254 222
rect 256 218 257 222
rect 256 214 261 218
rect 269 214 270 222
rect 272 214 275 222
rect 277 214 278 222
rect 295 214 296 222
rect 298 214 299 222
rect 311 214 312 222
rect 314 218 315 222
rect 314 214 319 218
rect 327 214 328 222
rect 330 214 333 222
rect 335 214 336 222
rect 348 214 349 222
rect 351 214 352 222
rect 364 214 365 222
rect 367 214 370 222
rect 372 214 373 222
rect 385 214 386 222
rect 388 218 389 222
rect 388 214 393 218
rect 401 214 402 222
rect 404 214 407 222
rect 409 214 410 222
rect 427 214 428 222
rect 430 214 431 222
rect 443 214 444 222
rect 446 218 447 222
rect 446 214 451 218
rect 459 214 460 222
rect 462 214 465 222
rect 467 214 468 222
rect 480 214 481 222
rect 483 214 484 222
<< ndcontact >>
rect 96 191 100 195
rect 109 191 113 195
rect 117 191 121 195
rect 125 191 129 195
rect 133 191 137 195
rect 146 191 150 195
rect 159 191 163 195
rect 167 191 171 195
rect 175 191 179 195
rect 183 191 187 195
rect 191 191 195 195
rect 204 191 208 195
rect 212 191 216 195
rect 220 191 224 195
rect 228 191 232 195
rect 241 191 245 195
rect 249 191 253 195
rect 257 191 261 195
rect 265 191 269 195
rect 278 191 282 195
rect 291 191 295 195
rect 299 191 303 195
rect 307 191 311 195
rect 315 191 319 195
rect 323 191 327 195
rect 336 191 340 195
rect 344 191 348 195
rect 352 191 356 195
rect 360 191 364 195
rect 373 191 377 195
rect 381 191 385 195
rect 389 191 393 195
rect 397 191 401 195
rect 410 191 414 195
rect 423 191 427 195
rect 431 191 435 195
rect 439 191 443 195
rect 447 191 451 195
rect 455 191 459 195
rect 468 191 472 195
rect 476 191 480 195
rect 484 191 488 195
<< pdcontact >>
rect 96 214 100 222
rect 109 214 113 222
rect 117 214 121 222
rect 125 218 129 222
rect 133 214 137 222
rect 146 214 150 222
rect 159 214 163 222
rect 167 214 171 222
rect 175 214 179 222
rect 183 218 187 222
rect 191 214 195 222
rect 204 214 208 222
rect 212 214 216 222
rect 220 214 224 222
rect 228 214 232 222
rect 241 214 245 222
rect 249 214 253 222
rect 257 218 261 222
rect 265 214 269 222
rect 278 214 282 222
rect 291 214 295 222
rect 299 214 303 222
rect 307 214 311 222
rect 315 218 319 222
rect 323 214 327 222
rect 336 214 340 222
rect 344 214 348 222
rect 352 214 356 222
rect 360 214 364 222
rect 373 214 377 222
rect 381 214 385 222
rect 389 218 393 222
rect 397 214 401 222
rect 410 214 414 222
rect 423 214 427 222
rect 431 214 435 222
rect 439 214 443 222
rect 447 218 451 222
rect 455 214 459 222
rect 468 214 472 222
rect 476 214 480 222
rect 484 214 488 222
<< psubstratepcontact >>
rect 126 175 130 179
rect 154 175 158 179
rect 184 175 188 179
rect 258 175 262 179
rect 286 175 290 179
rect 316 175 320 179
rect 390 175 394 179
rect 418 175 422 179
rect 448 175 452 179
<< nsubstratencontact >>
rect 126 232 130 236
rect 154 232 158 236
rect 184 232 188 236
rect 221 232 225 236
rect 258 232 262 236
rect 286 232 290 236
rect 316 232 320 236
rect 353 232 357 236
rect 390 232 394 236
rect 418 232 422 236
rect 448 232 452 236
rect 485 232 489 236
<< polysilicon >>
rect 101 222 103 224
rect 106 222 108 225
rect 122 222 124 224
rect 138 222 140 224
rect 143 222 145 225
rect 164 222 166 225
rect 180 222 182 225
rect 196 222 198 224
rect 201 222 203 225
rect 217 222 219 224
rect 233 222 235 224
rect 238 222 240 225
rect 254 222 256 224
rect 270 222 272 224
rect 275 222 277 225
rect 296 222 298 225
rect 312 222 314 225
rect 328 222 330 224
rect 333 222 335 225
rect 349 222 351 224
rect 365 222 367 224
rect 370 222 372 225
rect 386 222 388 224
rect 402 222 404 224
rect 407 222 409 225
rect 428 222 430 225
rect 444 222 446 225
rect 460 222 462 224
rect 465 222 467 225
rect 481 222 483 224
rect 101 209 103 214
rect 106 212 108 214
rect 101 195 103 205
rect 106 195 108 202
rect 122 195 124 214
rect 138 205 140 214
rect 143 212 145 214
rect 164 212 166 214
rect 180 211 182 214
rect 138 195 140 198
rect 143 195 145 197
rect 164 195 166 197
rect 180 195 182 207
rect 196 205 198 214
rect 201 212 203 214
rect 217 206 219 214
rect 233 209 235 214
rect 238 212 240 214
rect 196 195 198 198
rect 201 195 203 197
rect 217 195 219 202
rect 233 195 235 205
rect 238 195 240 202
rect 254 195 256 214
rect 270 205 272 214
rect 275 212 277 214
rect 296 212 298 214
rect 312 211 314 214
rect 270 195 272 198
rect 275 195 277 197
rect 296 195 298 197
rect 312 195 314 207
rect 328 205 330 214
rect 333 212 335 214
rect 349 206 351 214
rect 365 209 367 214
rect 370 212 372 214
rect 328 195 330 198
rect 333 195 335 197
rect 349 195 351 202
rect 365 195 367 205
rect 370 195 372 202
rect 386 195 388 214
rect 402 205 404 214
rect 407 212 409 214
rect 428 212 430 214
rect 444 211 446 214
rect 402 195 404 198
rect 407 195 409 197
rect 428 195 430 197
rect 444 195 446 207
rect 460 205 462 214
rect 465 212 467 214
rect 481 206 483 214
rect 460 195 462 198
rect 465 195 467 197
rect 481 195 483 202
rect 101 189 103 191
rect 106 188 108 191
rect 122 189 124 191
rect 138 189 140 191
rect 143 186 145 191
rect 164 186 166 191
rect 180 189 182 191
rect 196 189 198 191
rect 201 186 203 191
rect 217 189 219 191
rect 233 189 235 191
rect 238 188 240 191
rect 254 189 256 191
rect 270 189 272 191
rect 275 186 277 191
rect 296 186 298 191
rect 312 189 314 191
rect 328 189 330 191
rect 333 186 335 191
rect 349 189 351 191
rect 365 189 367 191
rect 370 188 372 191
rect 386 189 388 191
rect 402 189 404 191
rect 407 186 409 191
rect 428 186 430 191
rect 444 189 446 191
rect 460 189 462 191
rect 465 186 467 191
rect 481 189 483 191
<< polycontact >>
rect 106 225 110 229
rect 143 225 147 229
rect 163 225 167 229
rect 201 225 205 229
rect 238 225 242 229
rect 275 225 279 229
rect 295 225 299 229
rect 333 225 337 229
rect 370 225 374 229
rect 407 225 411 229
rect 427 225 431 229
rect 465 225 469 229
rect 100 205 104 209
rect 118 207 122 211
rect 178 207 182 211
rect 136 198 140 205
rect 194 198 198 205
rect 215 202 219 206
rect 232 205 236 209
rect 250 207 254 211
rect 310 207 314 211
rect 268 198 272 205
rect 326 198 330 205
rect 347 202 351 206
rect 364 205 368 209
rect 382 207 386 211
rect 442 207 446 211
rect 400 198 404 205
rect 458 198 462 205
rect 479 202 483 206
rect 106 184 110 188
rect 143 182 147 186
rect 163 182 167 186
rect 199 182 203 186
rect 238 184 242 188
rect 275 182 279 186
rect 295 182 299 186
rect 331 182 335 186
rect 370 184 374 188
rect 407 182 411 186
rect 427 182 431 186
rect 463 182 467 186
<< metal1 >>
rect 93 239 102 243
rect 106 239 138 243
rect 142 239 205 243
rect 209 239 234 243
rect 238 239 270 243
rect 274 239 337 243
rect 341 239 366 243
rect 370 239 402 243
rect 406 239 469 243
rect 473 239 489 243
rect 93 232 126 236
rect 130 232 154 236
rect 158 232 184 236
rect 188 232 221 236
rect 225 232 258 236
rect 262 232 286 236
rect 290 232 316 236
rect 320 232 353 236
rect 357 232 390 236
rect 394 232 418 236
rect 422 232 448 236
rect 452 232 485 236
rect 96 222 99 232
rect 117 222 120 232
rect 133 222 136 232
rect 147 225 152 229
rect 156 225 163 229
rect 175 222 178 232
rect 191 222 194 232
rect 212 222 215 232
rect 228 222 231 232
rect 249 222 252 232
rect 265 222 268 232
rect 279 225 284 229
rect 288 225 295 229
rect 307 222 310 232
rect 323 222 326 232
rect 344 222 347 232
rect 360 222 363 232
rect 381 222 384 232
rect 397 222 400 232
rect 411 225 416 229
rect 420 225 427 229
rect 439 222 442 232
rect 455 222 458 232
rect 476 222 479 232
rect 113 208 118 211
rect 122 208 146 211
rect 171 208 178 211
rect 182 208 204 211
rect 129 198 136 201
rect 140 202 159 205
rect 159 195 162 201
rect 187 198 194 201
rect 198 202 215 205
rect 245 208 250 211
rect 254 208 278 211
rect 303 208 310 211
rect 314 208 336 211
rect 261 198 268 201
rect 272 202 291 205
rect 291 195 294 201
rect 319 198 326 201
rect 330 202 347 205
rect 377 208 382 211
rect 386 208 410 211
rect 435 208 442 211
rect 446 208 468 211
rect 393 198 400 201
rect 404 202 423 205
rect 423 195 426 201
rect 451 198 458 201
rect 462 202 479 205
rect 96 179 99 191
rect 117 179 120 191
rect 133 179 136 191
rect 147 182 159 185
rect 175 179 178 191
rect 191 179 194 191
rect 212 179 215 191
rect 228 179 231 191
rect 249 179 252 191
rect 265 179 268 191
rect 279 182 291 185
rect 307 179 310 191
rect 323 179 326 191
rect 344 179 347 191
rect 360 179 363 191
rect 381 179 384 191
rect 397 179 400 191
rect 411 182 423 185
rect 439 179 442 191
rect 455 179 458 191
rect 476 179 479 191
rect 93 175 126 179
rect 130 175 154 179
rect 158 175 184 179
rect 188 175 258 179
rect 262 175 286 179
rect 290 175 316 179
rect 320 175 390 179
rect 394 175 418 179
rect 422 175 448 179
rect 452 175 489 179
rect 93 168 102 172
rect 106 168 153 172
rect 157 168 203 172
rect 207 168 234 172
rect 238 168 285 172
rect 289 168 335 172
rect 339 168 366 172
rect 370 168 417 172
rect 421 168 467 172
rect 471 168 489 172
<< m2contact >>
rect 102 239 106 243
rect 138 239 142 243
rect 205 239 209 243
rect 234 239 238 243
rect 270 239 274 243
rect 337 239 341 243
rect 366 239 370 243
rect 402 239 406 243
rect 469 239 473 243
rect 102 225 106 229
rect 152 225 156 229
rect 205 225 209 229
rect 234 225 238 229
rect 284 225 288 229
rect 337 225 341 229
rect 366 225 370 229
rect 416 225 420 229
rect 469 225 473 229
rect 125 214 129 218
rect 96 205 100 209
rect 109 208 113 214
rect 146 208 150 214
rect 159 210 163 214
rect 183 214 187 218
rect 257 214 261 218
rect 167 208 171 214
rect 204 208 208 214
rect 220 210 224 214
rect 109 195 113 199
rect 125 195 129 201
rect 159 201 163 205
rect 146 195 150 199
rect 167 195 171 199
rect 183 195 187 201
rect 228 205 232 209
rect 241 208 245 214
rect 278 208 282 214
rect 291 210 295 214
rect 315 214 319 218
rect 389 214 393 218
rect 299 208 303 214
rect 336 208 340 214
rect 352 210 356 214
rect 204 195 208 199
rect 220 195 224 199
rect 241 195 245 199
rect 257 195 261 201
rect 291 201 295 205
rect 278 195 282 199
rect 299 195 303 199
rect 315 195 319 201
rect 360 205 364 209
rect 373 208 377 214
rect 410 208 414 214
rect 423 210 427 214
rect 447 214 451 218
rect 431 208 435 214
rect 468 208 472 214
rect 484 210 488 214
rect 336 195 340 199
rect 352 195 356 199
rect 373 195 377 199
rect 389 195 393 201
rect 423 201 427 205
rect 410 195 414 199
rect 431 195 435 199
rect 447 195 451 201
rect 468 195 472 199
rect 484 195 488 199
rect 102 184 106 188
rect 139 182 143 186
rect 159 182 163 186
rect 203 182 207 186
rect 234 184 238 188
rect 271 182 275 186
rect 291 182 295 186
rect 335 182 339 186
rect 366 184 370 188
rect 403 182 407 186
rect 423 182 427 186
rect 467 182 471 186
rect 102 168 106 172
rect 153 168 157 172
rect 203 168 207 172
rect 234 168 238 172
rect 285 168 289 172
rect 335 168 339 172
rect 366 168 370 172
rect 417 168 421 172
rect 467 168 471 172
<< metal2 >>
rect 103 229 106 239
rect 93 205 96 208
rect 110 199 113 208
rect 126 201 129 214
rect 139 186 142 239
rect 206 229 209 239
rect 235 229 238 239
rect 146 214 150 218
rect 147 199 150 208
rect 102 172 105 184
rect 143 182 144 186
rect 153 172 156 225
rect 159 205 162 210
rect 168 199 171 208
rect 184 201 187 214
rect 205 199 208 208
rect 221 208 224 210
rect 221 205 228 208
rect 221 199 224 205
rect 242 199 245 208
rect 258 201 261 214
rect 204 172 207 182
rect 271 186 274 239
rect 338 229 341 239
rect 367 229 370 239
rect 278 214 282 218
rect 279 199 282 208
rect 234 172 237 184
rect 275 182 276 186
rect 285 172 288 225
rect 291 205 294 210
rect 300 199 303 208
rect 316 201 319 214
rect 337 199 340 208
rect 353 208 356 210
rect 353 205 360 208
rect 353 199 356 205
rect 374 199 377 208
rect 390 201 393 214
rect 336 172 339 182
rect 403 186 406 239
rect 470 229 473 239
rect 410 214 414 218
rect 411 199 414 208
rect 366 172 369 184
rect 407 182 408 186
rect 417 172 420 225
rect 423 205 426 210
rect 432 199 435 208
rect 448 201 451 214
rect 469 199 472 208
rect 485 208 488 210
rect 485 205 489 208
rect 485 199 488 205
rect 468 172 471 182
<< labels >>
rlabel metal1 96 232 99 236 1 Vdd!
rlabel metal1 97 175 100 179 1 GND!
rlabel metal1 98 168 101 172 2 ~clk
rlabel metal1 96 239 99 243 4 clk
rlabel metal2 94 207 94 207 3 D
rlabel metal2 223 207 223 207 1 q0
rlabel metal1 228 232 231 236 1 Vdd!
rlabel metal1 229 175 232 179 1 GND!
rlabel metal1 230 168 233 172 2 ~clk
rlabel metal1 228 239 231 243 4 clk
rlabel metal1 360 232 363 236 1 Vdd!
rlabel metal1 361 175 364 179 1 GND!
rlabel metal1 362 168 365 172 2 ~clk
rlabel metal1 360 239 363 243 4 clk
rlabel metal2 356 207 356 207 1 q1
rlabel metal2 486 207 486 207 7 q2
<< end >>
