magic
tech scmos
timestamp 1607474146
<< ntransistor >>
rect 50 144 52 148
rect 56 144 58 148
rect 72 144 74 148
rect 88 144 90 148
rect 94 144 96 148
rect 110 144 112 148
rect 131 144 133 148
rect 137 144 139 148
rect 153 144 155 148
rect 169 144 171 148
rect 175 144 177 148
rect 191 144 193 148
rect 109 120 111 124
rect 133 120 135 124
rect 129 109 131 113
rect 120 95 124 97
rect 109 86 111 90
rect 133 86 135 90
rect 218 31 220 35
rect 224 31 226 35
rect 240 31 242 35
rect 256 31 258 35
rect 262 31 264 35
rect 278 31 280 35
rect 299 31 301 35
rect 305 31 307 35
rect 321 31 323 35
rect 337 31 339 35
rect 343 31 345 35
rect 359 31 361 35
rect 50 12 52 16
rect 56 12 58 16
rect 72 12 74 16
rect 88 12 90 16
rect 94 12 96 16
rect 110 12 112 16
rect 131 12 133 16
rect 137 12 139 16
rect 153 12 155 16
rect 169 12 171 16
rect 175 12 177 16
rect 191 12 193 16
rect 277 7 279 11
rect 301 7 303 11
rect 297 -4 299 0
rect 50 -20 52 -16
rect 56 -20 58 -16
rect 72 -20 74 -16
rect 88 -20 90 -16
rect 94 -20 96 -16
rect 110 -20 112 -16
rect 131 -20 133 -16
rect 137 -20 139 -16
rect 153 -20 155 -16
rect 169 -20 171 -16
rect 175 -20 177 -16
rect 191 -20 193 -16
rect 288 -18 292 -16
rect 277 -27 279 -23
rect 301 -27 303 -23
rect 386 -82 388 -78
rect 392 -82 394 -78
rect 408 -82 410 -78
rect 424 -82 426 -78
rect 430 -82 432 -78
rect 446 -82 448 -78
rect 467 -82 469 -78
rect 473 -82 475 -78
rect 489 -82 491 -78
rect 505 -82 507 -78
rect 511 -82 513 -78
rect 527 -82 529 -78
rect 218 -101 220 -97
rect 224 -101 226 -97
rect 240 -101 242 -97
rect 256 -101 258 -97
rect 262 -101 264 -97
rect 278 -101 280 -97
rect 299 -101 301 -97
rect 305 -101 307 -97
rect 321 -101 323 -97
rect 337 -101 339 -97
rect 343 -101 345 -97
rect 359 -101 361 -97
rect 445 -106 447 -102
rect 469 -106 471 -102
rect 465 -117 467 -113
rect 218 -133 220 -129
rect 224 -133 226 -129
rect 240 -133 242 -129
rect 256 -133 258 -129
rect 262 -133 264 -129
rect 278 -133 280 -129
rect 299 -133 301 -129
rect 305 -133 307 -129
rect 321 -133 323 -129
rect 337 -133 339 -129
rect 343 -133 345 -129
rect 359 -133 361 -129
rect 456 -131 460 -129
rect 445 -140 447 -136
rect 469 -140 471 -136
rect 386 -214 388 -210
rect 392 -214 394 -210
rect 408 -214 410 -210
rect 424 -214 426 -210
rect 430 -214 432 -210
rect 446 -214 448 -210
rect 467 -214 469 -210
rect 473 -214 475 -210
rect 489 -214 491 -210
rect 505 -214 507 -210
rect 511 -214 513 -210
rect 527 -214 529 -210
rect 386 -230 388 -226
rect 392 -230 394 -226
rect 408 -230 410 -226
rect 424 -230 426 -226
rect 430 -230 432 -226
rect 446 -230 448 -226
rect 467 -230 469 -226
rect 473 -230 475 -226
rect 489 -230 491 -226
rect 505 -230 507 -226
rect 511 -230 513 -226
rect 527 -230 529 -226
<< ptransistor >>
rect 50 190 52 198
rect 56 190 58 198
rect 72 190 74 198
rect 88 190 90 198
rect 94 190 96 198
rect 110 190 112 198
rect 131 190 133 198
rect 137 190 139 198
rect 153 190 155 198
rect 169 190 171 198
rect 175 190 177 198
rect 191 190 193 198
rect 218 77 220 85
rect 224 77 226 85
rect 240 77 242 85
rect 256 77 258 85
rect 262 77 264 85
rect 278 77 280 85
rect 299 77 301 85
rect 305 77 307 85
rect 321 77 323 85
rect 337 77 339 85
rect 343 77 345 85
rect 359 77 361 85
rect 50 58 52 66
rect 56 58 58 66
rect 72 58 74 66
rect 88 58 90 66
rect 94 58 96 66
rect 110 58 112 66
rect 131 58 133 66
rect 137 58 139 66
rect 153 58 155 66
rect 169 58 171 66
rect 175 58 177 66
rect 191 58 193 66
rect 386 -36 388 -28
rect 392 -36 394 -28
rect 408 -36 410 -28
rect 424 -36 426 -28
rect 430 -36 432 -28
rect 446 -36 448 -28
rect 467 -36 469 -28
rect 473 -36 475 -28
rect 489 -36 491 -28
rect 505 -36 507 -28
rect 511 -36 513 -28
rect 527 -36 529 -28
rect 218 -55 220 -47
rect 224 -55 226 -47
rect 240 -55 242 -47
rect 256 -55 258 -47
rect 262 -55 264 -47
rect 278 -55 280 -47
rect 299 -55 301 -47
rect 305 -55 307 -47
rect 321 -55 323 -47
rect 337 -55 339 -47
rect 343 -55 345 -47
rect 359 -55 361 -47
rect 50 -70 52 -62
rect 56 -70 58 -62
rect 72 -70 74 -62
rect 88 -70 90 -62
rect 94 -70 96 -62
rect 110 -70 112 -62
rect 131 -70 133 -62
rect 137 -70 139 -62
rect 153 -70 155 -62
rect 169 -70 171 -62
rect 175 -70 177 -62
rect 191 -70 193 -62
rect 386 -168 388 -160
rect 392 -168 394 -160
rect 408 -168 410 -160
rect 424 -168 426 -160
rect 430 -168 432 -160
rect 446 -168 448 -160
rect 467 -168 469 -160
rect 473 -168 475 -160
rect 489 -168 491 -160
rect 505 -168 507 -160
rect 511 -168 513 -160
rect 527 -168 529 -160
rect 218 -183 220 -175
rect 224 -183 226 -175
rect 240 -183 242 -175
rect 256 -183 258 -175
rect 262 -183 264 -175
rect 278 -183 280 -175
rect 299 -183 301 -175
rect 305 -183 307 -175
rect 321 -183 323 -175
rect 337 -183 339 -175
rect 343 -183 345 -175
rect 359 -183 361 -175
rect 386 -280 388 -272
rect 392 -280 394 -272
rect 408 -280 410 -272
rect 424 -280 426 -272
rect 430 -280 432 -272
rect 446 -280 448 -272
rect 467 -280 469 -272
rect 473 -280 475 -272
rect 489 -280 491 -272
rect 505 -280 507 -272
rect 511 -280 513 -272
rect 527 -280 529 -272
<< ndiffusion >>
rect 49 144 50 148
rect 52 144 56 148
rect 58 144 59 148
rect 71 144 72 148
rect 74 144 75 148
rect 87 144 88 148
rect 90 144 94 148
rect 96 144 97 148
rect 109 144 110 148
rect 112 144 113 148
rect 130 144 131 148
rect 133 144 137 148
rect 139 144 140 148
rect 152 144 153 148
rect 155 144 156 148
rect 168 144 169 148
rect 171 144 175 148
rect 177 144 178 148
rect 190 144 191 148
rect 193 144 194 148
rect 108 120 109 124
rect 111 120 112 124
rect 132 120 133 124
rect 135 120 136 124
rect 128 109 129 113
rect 131 109 132 113
rect 120 97 124 98
rect 120 94 124 95
rect 108 86 109 90
rect 111 86 112 90
rect 132 86 133 90
rect 135 86 136 90
rect 217 31 218 35
rect 220 31 224 35
rect 226 31 227 35
rect 239 31 240 35
rect 242 31 243 35
rect 255 31 256 35
rect 258 31 262 35
rect 264 31 265 35
rect 277 31 278 35
rect 280 31 281 35
rect 298 31 299 35
rect 301 31 305 35
rect 307 31 308 35
rect 320 31 321 35
rect 323 31 324 35
rect 336 31 337 35
rect 339 31 343 35
rect 345 31 346 35
rect 358 31 359 35
rect 361 31 362 35
rect 49 12 50 16
rect 52 12 56 16
rect 58 12 59 16
rect 71 12 72 16
rect 74 12 75 16
rect 87 12 88 16
rect 90 12 94 16
rect 96 12 97 16
rect 109 12 110 16
rect 112 12 113 16
rect 130 12 131 16
rect 133 12 137 16
rect 139 12 140 16
rect 152 12 153 16
rect 155 12 156 16
rect 168 12 169 16
rect 171 12 175 16
rect 177 12 178 16
rect 190 12 191 16
rect 193 12 194 16
rect 276 7 277 11
rect 279 7 280 11
rect 300 7 301 11
rect 303 7 304 11
rect 296 -4 297 0
rect 299 -4 300 0
rect 49 -20 50 -16
rect 52 -20 56 -16
rect 58 -20 59 -16
rect 71 -20 72 -16
rect 74 -20 75 -16
rect 87 -20 88 -16
rect 90 -20 94 -16
rect 96 -20 97 -16
rect 109 -20 110 -16
rect 112 -20 113 -16
rect 130 -20 131 -16
rect 133 -20 137 -16
rect 139 -20 140 -16
rect 152 -20 153 -16
rect 155 -20 156 -16
rect 168 -20 169 -16
rect 171 -20 175 -16
rect 177 -20 178 -16
rect 190 -20 191 -16
rect 193 -20 194 -16
rect 288 -16 292 -15
rect 288 -19 292 -18
rect 276 -27 277 -23
rect 279 -27 280 -23
rect 300 -27 301 -23
rect 303 -27 304 -23
rect 385 -82 386 -78
rect 388 -82 392 -78
rect 394 -82 395 -78
rect 407 -82 408 -78
rect 410 -82 411 -78
rect 423 -82 424 -78
rect 426 -82 430 -78
rect 432 -82 433 -78
rect 445 -82 446 -78
rect 448 -82 449 -78
rect 466 -82 467 -78
rect 469 -82 473 -78
rect 475 -82 476 -78
rect 488 -82 489 -78
rect 491 -82 492 -78
rect 504 -82 505 -78
rect 507 -82 511 -78
rect 513 -82 514 -78
rect 526 -82 527 -78
rect 529 -82 530 -78
rect 217 -101 218 -97
rect 220 -101 224 -97
rect 226 -101 227 -97
rect 239 -101 240 -97
rect 242 -101 243 -97
rect 255 -101 256 -97
rect 258 -101 262 -97
rect 264 -101 265 -97
rect 277 -101 278 -97
rect 280 -101 281 -97
rect 298 -101 299 -97
rect 301 -101 305 -97
rect 307 -101 308 -97
rect 320 -101 321 -97
rect 323 -101 324 -97
rect 336 -101 337 -97
rect 339 -101 343 -97
rect 345 -101 346 -97
rect 358 -101 359 -97
rect 361 -101 362 -97
rect 444 -106 445 -102
rect 447 -106 448 -102
rect 468 -106 469 -102
rect 471 -106 472 -102
rect 464 -117 465 -113
rect 467 -117 468 -113
rect 217 -133 218 -129
rect 220 -133 224 -129
rect 226 -133 227 -129
rect 239 -133 240 -129
rect 242 -133 243 -129
rect 255 -133 256 -129
rect 258 -133 262 -129
rect 264 -133 265 -129
rect 277 -133 278 -129
rect 280 -133 281 -129
rect 298 -133 299 -129
rect 301 -133 305 -129
rect 307 -133 308 -129
rect 320 -133 321 -129
rect 323 -133 324 -129
rect 336 -133 337 -129
rect 339 -133 343 -129
rect 345 -133 346 -129
rect 358 -133 359 -129
rect 361 -133 362 -129
rect 456 -129 460 -128
rect 456 -132 460 -131
rect 444 -140 445 -136
rect 447 -140 448 -136
rect 468 -140 469 -136
rect 471 -140 472 -136
rect 385 -214 386 -210
rect 388 -214 392 -210
rect 394 -214 395 -210
rect 407 -214 408 -210
rect 410 -214 411 -210
rect 423 -214 424 -210
rect 426 -214 430 -210
rect 432 -214 433 -210
rect 445 -214 446 -210
rect 448 -214 449 -210
rect 466 -214 467 -210
rect 469 -214 473 -210
rect 475 -214 476 -210
rect 488 -214 489 -210
rect 491 -214 492 -210
rect 504 -214 505 -210
rect 507 -214 511 -210
rect 513 -214 514 -210
rect 526 -214 527 -210
rect 529 -214 530 -210
rect 385 -230 386 -226
rect 388 -230 392 -226
rect 394 -230 395 -226
rect 407 -230 408 -226
rect 410 -230 411 -226
rect 423 -230 424 -226
rect 426 -230 430 -226
rect 432 -230 433 -226
rect 445 -230 446 -226
rect 448 -230 449 -226
rect 466 -230 467 -226
rect 469 -230 473 -226
rect 475 -230 476 -226
rect 488 -230 489 -226
rect 491 -230 492 -226
rect 504 -230 505 -226
rect 507 -230 511 -226
rect 513 -230 514 -226
rect 526 -230 527 -226
rect 529 -230 530 -226
<< pdiffusion >>
rect 49 190 50 198
rect 52 190 56 198
rect 58 194 59 198
rect 58 190 63 194
rect 71 190 72 198
rect 74 194 75 198
rect 74 190 79 194
rect 87 190 88 198
rect 90 190 94 198
rect 96 194 97 198
rect 96 190 101 194
rect 109 190 110 198
rect 112 194 113 198
rect 112 190 117 194
rect 130 190 131 198
rect 133 190 137 198
rect 139 194 140 198
rect 139 190 144 194
rect 152 190 153 198
rect 155 194 156 198
rect 155 190 160 194
rect 168 190 169 198
rect 171 190 175 198
rect 177 194 178 198
rect 177 190 182 194
rect 190 190 191 198
rect 193 194 194 198
rect 193 190 198 194
rect 217 77 218 85
rect 220 77 224 85
rect 226 81 227 85
rect 226 77 231 81
rect 239 77 240 85
rect 242 81 243 85
rect 242 77 247 81
rect 255 77 256 85
rect 258 77 262 85
rect 264 81 265 85
rect 264 77 269 81
rect 277 77 278 85
rect 280 81 281 85
rect 280 77 285 81
rect 298 77 299 85
rect 301 77 305 85
rect 307 81 308 85
rect 307 77 312 81
rect 320 77 321 85
rect 323 81 324 85
rect 323 77 328 81
rect 336 77 337 85
rect 339 77 343 85
rect 345 81 346 85
rect 345 77 350 81
rect 358 77 359 85
rect 361 81 362 85
rect 361 77 366 81
rect 49 58 50 66
rect 52 58 56 66
rect 58 62 59 66
rect 58 58 63 62
rect 71 58 72 66
rect 74 62 75 66
rect 74 58 79 62
rect 87 58 88 66
rect 90 58 94 66
rect 96 62 97 66
rect 96 58 101 62
rect 109 58 110 66
rect 112 62 113 66
rect 112 58 117 62
rect 130 58 131 66
rect 133 58 137 66
rect 139 62 140 66
rect 139 58 144 62
rect 152 58 153 66
rect 155 62 156 66
rect 155 58 160 62
rect 168 58 169 66
rect 171 58 175 66
rect 177 62 178 66
rect 177 58 182 62
rect 190 58 191 66
rect 193 62 194 66
rect 193 58 198 62
rect 385 -36 386 -28
rect 388 -36 392 -28
rect 394 -32 395 -28
rect 394 -36 399 -32
rect 407 -36 408 -28
rect 410 -32 411 -28
rect 410 -36 415 -32
rect 423 -36 424 -28
rect 426 -36 430 -28
rect 432 -32 433 -28
rect 432 -36 437 -32
rect 445 -36 446 -28
rect 448 -32 449 -28
rect 448 -36 453 -32
rect 466 -36 467 -28
rect 469 -36 473 -28
rect 475 -32 476 -28
rect 475 -36 480 -32
rect 488 -36 489 -28
rect 491 -32 492 -28
rect 491 -36 496 -32
rect 504 -36 505 -28
rect 507 -36 511 -28
rect 513 -32 514 -28
rect 513 -36 518 -32
rect 526 -36 527 -28
rect 529 -32 530 -28
rect 529 -36 534 -32
rect 217 -55 218 -47
rect 220 -55 224 -47
rect 226 -51 227 -47
rect 226 -55 231 -51
rect 239 -55 240 -47
rect 242 -51 243 -47
rect 242 -55 247 -51
rect 255 -55 256 -47
rect 258 -55 262 -47
rect 264 -51 265 -47
rect 264 -55 269 -51
rect 277 -55 278 -47
rect 280 -51 281 -47
rect 280 -55 285 -51
rect 298 -55 299 -47
rect 301 -55 305 -47
rect 307 -51 308 -47
rect 307 -55 312 -51
rect 320 -55 321 -47
rect 323 -51 324 -47
rect 323 -55 328 -51
rect 336 -55 337 -47
rect 339 -55 343 -47
rect 345 -51 346 -47
rect 345 -55 350 -51
rect 358 -55 359 -47
rect 361 -51 362 -47
rect 361 -55 366 -51
rect 49 -70 50 -62
rect 52 -70 56 -62
rect 58 -66 63 -62
rect 58 -70 59 -66
rect 71 -70 72 -62
rect 74 -66 79 -62
rect 74 -70 75 -66
rect 87 -70 88 -62
rect 90 -70 94 -62
rect 96 -66 101 -62
rect 96 -70 97 -66
rect 109 -70 110 -62
rect 112 -66 117 -62
rect 112 -70 113 -66
rect 130 -70 131 -62
rect 133 -70 137 -62
rect 139 -66 144 -62
rect 139 -70 140 -66
rect 152 -70 153 -62
rect 155 -66 160 -62
rect 155 -70 156 -66
rect 168 -70 169 -62
rect 171 -70 175 -62
rect 177 -66 182 -62
rect 177 -70 178 -66
rect 190 -70 191 -62
rect 193 -66 198 -62
rect 193 -70 194 -66
rect 385 -168 386 -160
rect 388 -168 392 -160
rect 394 -164 395 -160
rect 394 -168 399 -164
rect 407 -168 408 -160
rect 410 -164 411 -160
rect 410 -168 415 -164
rect 423 -168 424 -160
rect 426 -168 430 -160
rect 432 -164 433 -160
rect 432 -168 437 -164
rect 445 -168 446 -160
rect 448 -164 449 -160
rect 448 -168 453 -164
rect 466 -168 467 -160
rect 469 -168 473 -160
rect 475 -164 476 -160
rect 475 -168 480 -164
rect 488 -168 489 -160
rect 491 -164 492 -160
rect 491 -168 496 -164
rect 504 -168 505 -160
rect 507 -168 511 -160
rect 513 -164 514 -160
rect 513 -168 518 -164
rect 526 -168 527 -160
rect 529 -164 530 -160
rect 529 -168 534 -164
rect 217 -183 218 -175
rect 220 -183 224 -175
rect 226 -179 231 -175
rect 226 -183 227 -179
rect 239 -183 240 -175
rect 242 -179 247 -175
rect 242 -183 243 -179
rect 255 -183 256 -175
rect 258 -183 262 -175
rect 264 -179 269 -175
rect 264 -183 265 -179
rect 277 -183 278 -175
rect 280 -179 285 -175
rect 280 -183 281 -179
rect 298 -183 299 -175
rect 301 -183 305 -175
rect 307 -179 312 -175
rect 307 -183 308 -179
rect 320 -183 321 -175
rect 323 -179 328 -175
rect 323 -183 324 -179
rect 336 -183 337 -175
rect 339 -183 343 -175
rect 345 -179 350 -175
rect 345 -183 346 -179
rect 358 -183 359 -175
rect 361 -179 366 -175
rect 361 -183 362 -179
rect 385 -280 386 -272
rect 388 -280 392 -272
rect 394 -276 399 -272
rect 394 -280 395 -276
rect 407 -280 408 -272
rect 410 -276 415 -272
rect 410 -280 411 -276
rect 423 -280 424 -272
rect 426 -280 430 -272
rect 432 -276 437 -272
rect 432 -280 433 -276
rect 445 -280 446 -272
rect 448 -276 453 -272
rect 448 -280 449 -276
rect 466 -280 467 -272
rect 469 -280 473 -272
rect 475 -276 480 -272
rect 475 -280 476 -276
rect 488 -280 489 -272
rect 491 -276 496 -272
rect 491 -280 492 -276
rect 504 -280 505 -272
rect 507 -280 511 -272
rect 513 -276 518 -272
rect 513 -280 514 -276
rect 526 -280 527 -272
rect 529 -276 534 -272
rect 529 -280 530 -276
<< ndcontact >>
rect 45 144 49 148
rect 59 144 63 148
rect 67 144 71 148
rect 75 144 79 148
rect 83 144 87 148
rect 97 144 101 148
rect 105 144 109 148
rect 113 144 117 148
rect 126 144 130 148
rect 140 144 144 148
rect 148 144 152 148
rect 156 144 160 148
rect 164 144 168 148
rect 178 144 182 148
rect 186 144 190 148
rect 194 144 198 148
rect 104 120 108 124
rect 112 120 116 124
rect 128 120 132 124
rect 136 120 140 124
rect 124 109 128 113
rect 132 109 136 113
rect 120 98 124 102
rect 120 90 124 94
rect 104 86 108 90
rect 112 86 116 90
rect 128 86 132 90
rect 136 86 140 90
rect 213 31 217 35
rect 227 31 231 35
rect 235 31 239 35
rect 243 31 247 35
rect 251 31 255 35
rect 265 31 269 35
rect 273 31 277 35
rect 281 31 285 35
rect 294 31 298 35
rect 308 31 312 35
rect 316 31 320 35
rect 324 31 328 35
rect 332 31 336 35
rect 346 31 350 35
rect 354 31 358 35
rect 362 31 366 35
rect 45 12 49 16
rect 59 12 63 16
rect 67 12 71 16
rect 75 12 79 16
rect 83 12 87 16
rect 97 12 101 16
rect 105 12 109 16
rect 113 12 117 16
rect 126 12 130 16
rect 140 12 144 16
rect 148 12 152 16
rect 156 12 160 16
rect 164 12 168 16
rect 178 12 182 16
rect 186 12 190 16
rect 194 12 198 16
rect 272 7 276 11
rect 280 7 284 11
rect 296 7 300 11
rect 304 7 308 11
rect 292 -4 296 0
rect 300 -4 304 0
rect 45 -20 49 -16
rect 59 -20 63 -16
rect 67 -20 71 -16
rect 75 -20 79 -16
rect 83 -20 87 -16
rect 97 -20 101 -16
rect 105 -20 109 -16
rect 113 -20 117 -16
rect 126 -20 130 -16
rect 140 -20 144 -16
rect 148 -20 152 -16
rect 156 -20 160 -16
rect 164 -20 168 -16
rect 178 -20 182 -16
rect 186 -20 190 -16
rect 194 -20 198 -16
rect 288 -15 292 -11
rect 288 -23 292 -19
rect 272 -27 276 -23
rect 280 -27 284 -23
rect 296 -27 300 -23
rect 304 -27 308 -23
rect 381 -82 385 -78
rect 395 -82 399 -78
rect 403 -82 407 -78
rect 411 -82 415 -78
rect 419 -82 423 -78
rect 433 -82 437 -78
rect 441 -82 445 -78
rect 449 -82 453 -78
rect 462 -82 466 -78
rect 476 -82 480 -78
rect 484 -82 488 -78
rect 492 -82 496 -78
rect 500 -82 504 -78
rect 514 -82 518 -78
rect 522 -82 526 -78
rect 530 -82 534 -78
rect 213 -101 217 -97
rect 227 -101 231 -97
rect 235 -101 239 -97
rect 243 -101 247 -97
rect 251 -101 255 -97
rect 265 -101 269 -97
rect 273 -101 277 -97
rect 281 -101 285 -97
rect 294 -101 298 -97
rect 308 -101 312 -97
rect 316 -101 320 -97
rect 324 -101 328 -97
rect 332 -101 336 -97
rect 346 -101 350 -97
rect 354 -101 358 -97
rect 362 -101 366 -97
rect 440 -106 444 -102
rect 448 -106 452 -102
rect 464 -106 468 -102
rect 472 -106 476 -102
rect 460 -117 464 -113
rect 468 -117 472 -113
rect 213 -133 217 -129
rect 227 -133 231 -129
rect 235 -133 239 -129
rect 243 -133 247 -129
rect 251 -133 255 -129
rect 265 -133 269 -129
rect 273 -133 277 -129
rect 281 -133 285 -129
rect 294 -133 298 -129
rect 308 -133 312 -129
rect 316 -133 320 -129
rect 324 -133 328 -129
rect 332 -133 336 -129
rect 346 -133 350 -129
rect 354 -133 358 -129
rect 362 -133 366 -129
rect 456 -128 460 -124
rect 456 -136 460 -132
rect 440 -140 444 -136
rect 448 -140 452 -136
rect 464 -140 468 -136
rect 472 -140 476 -136
rect 381 -214 385 -210
rect 395 -214 399 -210
rect 403 -214 407 -210
rect 411 -214 415 -210
rect 419 -214 423 -210
rect 433 -214 437 -210
rect 441 -214 445 -210
rect 449 -214 453 -210
rect 462 -214 466 -210
rect 476 -214 480 -210
rect 484 -214 488 -210
rect 492 -214 496 -210
rect 500 -214 504 -210
rect 514 -214 518 -210
rect 522 -214 526 -210
rect 530 -214 534 -210
rect 381 -230 385 -226
rect 395 -230 399 -226
rect 403 -230 407 -226
rect 411 -230 415 -226
rect 419 -230 423 -226
rect 433 -230 437 -226
rect 441 -230 445 -226
rect 449 -230 453 -226
rect 462 -230 466 -226
rect 476 -230 480 -226
rect 484 -230 488 -226
rect 492 -230 496 -226
rect 500 -230 504 -226
rect 514 -230 518 -226
rect 522 -230 526 -226
rect 530 -230 534 -226
<< pdcontact >>
rect 45 190 49 198
rect 59 194 63 198
rect 67 190 71 198
rect 75 194 79 198
rect 83 190 87 198
rect 97 194 101 198
rect 105 190 109 198
rect 113 194 117 198
rect 126 190 130 198
rect 140 194 144 198
rect 148 190 152 198
rect 156 194 160 198
rect 164 190 168 198
rect 178 194 182 198
rect 186 190 190 198
rect 194 194 198 198
rect 213 77 217 85
rect 227 81 231 85
rect 235 77 239 85
rect 243 81 247 85
rect 251 77 255 85
rect 265 81 269 85
rect 273 77 277 85
rect 281 81 285 85
rect 294 77 298 85
rect 308 81 312 85
rect 316 77 320 85
rect 324 81 328 85
rect 332 77 336 85
rect 346 81 350 85
rect 354 77 358 85
rect 362 81 366 85
rect 45 58 49 66
rect 59 62 63 66
rect 67 58 71 66
rect 75 62 79 66
rect 83 58 87 66
rect 97 62 101 66
rect 105 58 109 66
rect 113 62 117 66
rect 126 58 130 66
rect 140 62 144 66
rect 148 58 152 66
rect 156 62 160 66
rect 164 58 168 66
rect 178 62 182 66
rect 186 58 190 66
rect 194 62 198 66
rect 381 -36 385 -28
rect 395 -32 399 -28
rect 403 -36 407 -28
rect 411 -32 415 -28
rect 419 -36 423 -28
rect 433 -32 437 -28
rect 441 -36 445 -28
rect 449 -32 453 -28
rect 462 -36 466 -28
rect 476 -32 480 -28
rect 484 -36 488 -28
rect 492 -32 496 -28
rect 500 -36 504 -28
rect 514 -32 518 -28
rect 522 -36 526 -28
rect 530 -32 534 -28
rect 213 -55 217 -47
rect 227 -51 231 -47
rect 235 -55 239 -47
rect 243 -51 247 -47
rect 251 -55 255 -47
rect 265 -51 269 -47
rect 273 -55 277 -47
rect 281 -51 285 -47
rect 294 -55 298 -47
rect 308 -51 312 -47
rect 316 -55 320 -47
rect 324 -51 328 -47
rect 332 -55 336 -47
rect 346 -51 350 -47
rect 354 -55 358 -47
rect 362 -51 366 -47
rect 45 -70 49 -62
rect 59 -70 63 -66
rect 67 -70 71 -62
rect 75 -70 79 -66
rect 83 -70 87 -62
rect 97 -70 101 -66
rect 105 -70 109 -62
rect 113 -70 117 -66
rect 126 -70 130 -62
rect 140 -70 144 -66
rect 148 -70 152 -62
rect 156 -70 160 -66
rect 164 -70 168 -62
rect 178 -70 182 -66
rect 186 -70 190 -62
rect 194 -70 198 -66
rect 381 -168 385 -160
rect 395 -164 399 -160
rect 403 -168 407 -160
rect 411 -164 415 -160
rect 419 -168 423 -160
rect 433 -164 437 -160
rect 441 -168 445 -160
rect 449 -164 453 -160
rect 462 -168 466 -160
rect 476 -164 480 -160
rect 484 -168 488 -160
rect 492 -164 496 -160
rect 500 -168 504 -160
rect 514 -164 518 -160
rect 522 -168 526 -160
rect 530 -164 534 -160
rect 213 -183 217 -175
rect 227 -183 231 -179
rect 235 -183 239 -175
rect 243 -183 247 -179
rect 251 -183 255 -175
rect 265 -183 269 -179
rect 273 -183 277 -175
rect 281 -183 285 -179
rect 294 -183 298 -175
rect 308 -183 312 -179
rect 316 -183 320 -175
rect 324 -183 328 -179
rect 332 -183 336 -175
rect 346 -183 350 -179
rect 354 -183 358 -175
rect 362 -183 366 -179
rect 381 -280 385 -272
rect 395 -280 399 -276
rect 403 -280 407 -272
rect 411 -280 415 -276
rect 419 -280 423 -272
rect 433 -280 437 -276
rect 441 -280 445 -272
rect 449 -280 453 -276
rect 462 -280 466 -272
rect 476 -280 480 -276
rect 484 -280 488 -272
rect 492 -280 496 -276
rect 500 -280 504 -272
rect 514 -280 518 -276
rect 522 -280 526 -272
rect 530 -280 534 -276
<< psubstratepcontact >>
rect 38 136 42 140
rect 80 136 84 140
rect 89 136 93 140
rect 101 136 105 140
rect 161 136 165 140
rect 170 136 174 140
rect 182 136 186 140
rect 206 23 210 27
rect 248 23 252 27
rect 257 23 261 27
rect 269 23 273 27
rect 329 23 333 27
rect 338 23 342 27
rect 350 23 354 27
rect 112 4 116 8
rect 143 4 147 8
rect 38 -12 42 -8
rect 80 -12 84 -8
rect 89 -12 93 -8
rect 101 -12 105 -8
rect 161 -12 165 -8
rect 170 -12 174 -8
rect 182 -12 186 -8
rect 374 -90 378 -86
rect 416 -90 420 -86
rect 425 -90 429 -86
rect 437 -90 441 -86
rect 497 -90 501 -86
rect 506 -90 510 -86
rect 518 -90 522 -86
rect 280 -109 284 -105
rect 311 -109 315 -105
rect 206 -125 210 -121
rect 248 -125 252 -121
rect 257 -125 261 -121
rect 269 -125 273 -121
rect 329 -125 333 -121
rect 338 -125 342 -121
rect 350 -125 354 -121
rect 374 -222 378 -218
rect 416 -222 420 -218
rect 425 -222 429 -218
rect 437 -222 441 -218
rect 448 -222 452 -218
rect 479 -222 483 -218
rect 497 -222 501 -218
rect 506 -222 510 -218
rect 518 -222 522 -218
<< nsubstratencontact >>
rect 45 202 49 206
rect 61 202 65 206
rect 76 202 80 206
rect 98 202 102 206
rect 126 202 130 206
rect 142 202 146 206
rect 157 202 161 206
rect 179 202 183 206
rect 213 89 217 93
rect 229 89 233 93
rect 244 89 248 93
rect 266 89 270 93
rect 294 89 298 93
rect 310 89 314 93
rect 325 89 329 93
rect 347 89 351 93
rect 45 70 49 74
rect 61 70 65 74
rect 76 70 80 74
rect 126 70 130 74
rect 142 70 146 74
rect 157 70 161 74
rect 179 70 183 74
rect 381 -24 385 -20
rect 397 -24 401 -20
rect 412 -24 416 -20
rect 434 -24 438 -20
rect 462 -24 466 -20
rect 478 -24 482 -20
rect 493 -24 497 -20
rect 515 -24 519 -20
rect 213 -43 217 -39
rect 229 -43 233 -39
rect 244 -43 248 -39
rect 294 -43 298 -39
rect 310 -43 314 -39
rect 325 -43 329 -39
rect 347 -43 351 -39
rect 45 -78 49 -74
rect 61 -78 65 -74
rect 76 -78 80 -74
rect 126 -78 130 -74
rect 142 -78 146 -74
rect 157 -78 161 -74
rect 179 -78 183 -74
rect 381 -156 385 -152
rect 397 -156 401 -152
rect 412 -156 416 -152
rect 462 -156 466 -152
rect 478 -156 482 -152
rect 493 -156 497 -152
rect 515 -156 519 -152
rect 213 -191 217 -187
rect 229 -191 233 -187
rect 244 -191 248 -187
rect 294 -191 298 -187
rect 310 -191 314 -187
rect 325 -191 329 -187
rect 347 -191 351 -187
rect 381 -288 385 -284
rect 397 -288 401 -284
rect 412 -288 416 -284
rect 462 -288 466 -284
rect 478 -288 482 -284
rect 493 -288 497 -284
rect 515 -288 519 -284
<< polysilicon >>
rect 50 198 52 200
rect 56 198 58 200
rect 72 198 74 200
rect 88 198 90 200
rect 94 198 96 200
rect 110 198 112 200
rect 131 198 133 200
rect 137 198 139 200
rect 153 198 155 200
rect 169 198 171 200
rect 175 198 177 200
rect 191 198 193 200
rect 50 173 52 190
rect 56 187 58 190
rect 72 173 74 190
rect 88 187 90 190
rect 50 148 52 169
rect 56 148 58 155
rect 72 148 74 169
rect 88 148 90 183
rect 94 180 96 190
rect 110 173 112 190
rect 131 173 133 190
rect 137 187 139 190
rect 153 173 155 190
rect 169 187 171 190
rect 94 148 96 162
rect 110 148 112 169
rect 131 148 133 169
rect 137 148 139 155
rect 153 148 155 169
rect 169 148 171 183
rect 175 180 177 190
rect 191 173 193 190
rect 175 148 177 162
rect 191 148 193 169
rect 50 142 52 144
rect 56 142 58 144
rect 72 142 74 144
rect 88 142 90 144
rect 94 142 96 144
rect 110 142 112 144
rect 131 142 133 144
rect 137 142 139 144
rect 153 142 155 144
rect 169 142 171 144
rect 175 142 177 144
rect 191 142 193 144
rect 109 124 111 128
rect 133 124 135 128
rect 109 118 111 120
rect 133 118 135 120
rect 129 113 131 115
rect 129 106 131 109
rect 117 96 120 97
rect 113 95 120 96
rect 124 95 126 97
rect 109 90 111 92
rect 133 90 135 92
rect 109 82 111 86
rect 133 82 135 86
rect 218 85 220 87
rect 224 85 226 87
rect 240 85 242 87
rect 256 85 258 87
rect 262 85 264 87
rect 278 85 280 87
rect 299 85 301 87
rect 305 85 307 87
rect 321 85 323 87
rect 337 85 339 87
rect 343 85 345 87
rect 359 85 361 87
rect 50 66 52 68
rect 56 66 58 68
rect 72 66 74 68
rect 88 66 90 68
rect 94 66 96 68
rect 110 66 112 68
rect 131 66 133 68
rect 137 66 139 68
rect 153 66 155 68
rect 169 66 171 68
rect 175 66 177 68
rect 191 66 193 68
rect 218 60 220 77
rect 224 74 226 77
rect 240 60 242 77
rect 256 74 258 77
rect 50 41 52 58
rect 56 55 58 58
rect 72 41 74 58
rect 88 55 90 58
rect 50 16 52 37
rect 56 16 58 23
rect 72 16 74 37
rect 88 16 90 51
rect 94 48 96 58
rect 110 41 112 58
rect 131 41 133 58
rect 137 55 139 58
rect 153 41 155 58
rect 169 55 171 58
rect 94 16 96 30
rect 110 16 112 37
rect 131 16 133 37
rect 137 16 139 23
rect 153 16 155 37
rect 169 16 171 51
rect 175 48 177 58
rect 191 41 193 58
rect 175 16 177 30
rect 191 16 193 37
rect 218 35 220 56
rect 224 35 226 42
rect 240 35 242 56
rect 256 35 258 70
rect 262 67 264 77
rect 278 60 280 77
rect 299 60 301 77
rect 305 74 307 77
rect 321 60 323 77
rect 337 74 339 77
rect 262 35 264 49
rect 278 35 280 56
rect 299 35 301 56
rect 305 35 307 42
rect 321 35 323 56
rect 337 35 339 70
rect 343 67 345 77
rect 359 60 361 77
rect 343 35 345 49
rect 359 35 361 56
rect 218 29 220 31
rect 224 29 226 31
rect 240 29 242 31
rect 256 29 258 31
rect 262 29 264 31
rect 278 29 280 31
rect 299 29 301 31
rect 305 29 307 31
rect 321 29 323 31
rect 337 29 339 31
rect 343 29 345 31
rect 359 29 361 31
rect 50 10 52 12
rect 56 10 58 12
rect 72 10 74 12
rect 88 10 90 12
rect 94 10 96 12
rect 110 10 112 12
rect 131 10 133 12
rect 137 10 139 12
rect 153 10 155 12
rect 169 10 171 12
rect 175 10 177 12
rect 191 10 193 12
rect 277 11 279 15
rect 301 11 303 15
rect 277 5 279 7
rect 301 5 303 7
rect 297 0 299 2
rect 297 -7 299 -4
rect 50 -16 52 -14
rect 56 -16 58 -14
rect 72 -16 74 -14
rect 88 -16 90 -14
rect 94 -16 96 -14
rect 110 -16 112 -14
rect 131 -16 133 -14
rect 137 -16 139 -14
rect 153 -16 155 -14
rect 169 -16 171 -14
rect 175 -16 177 -14
rect 191 -16 193 -14
rect 285 -17 288 -16
rect 281 -18 288 -17
rect 292 -18 294 -16
rect 50 -41 52 -20
rect 56 -27 58 -20
rect 72 -41 74 -20
rect 50 -62 52 -45
rect 56 -62 58 -59
rect 72 -62 74 -45
rect 88 -55 90 -20
rect 94 -34 96 -20
rect 110 -41 112 -20
rect 131 -41 133 -20
rect 137 -27 139 -20
rect 153 -41 155 -20
rect 88 -62 90 -59
rect 94 -62 96 -52
rect 110 -62 112 -45
rect 131 -62 133 -45
rect 137 -62 139 -59
rect 153 -62 155 -45
rect 169 -55 171 -20
rect 175 -34 177 -20
rect 191 -41 193 -20
rect 277 -23 279 -21
rect 301 -23 303 -21
rect 277 -31 279 -27
rect 301 -31 303 -27
rect 386 -28 388 -26
rect 392 -28 394 -26
rect 408 -28 410 -26
rect 424 -28 426 -26
rect 430 -28 432 -26
rect 446 -28 448 -26
rect 467 -28 469 -26
rect 473 -28 475 -26
rect 489 -28 491 -26
rect 505 -28 507 -26
rect 511 -28 513 -26
rect 527 -28 529 -26
rect 169 -62 171 -59
rect 175 -62 177 -52
rect 191 -62 193 -45
rect 218 -47 220 -45
rect 224 -47 226 -45
rect 240 -47 242 -45
rect 256 -47 258 -45
rect 262 -47 264 -45
rect 278 -47 280 -45
rect 299 -47 301 -45
rect 305 -47 307 -45
rect 321 -47 323 -45
rect 337 -47 339 -45
rect 343 -47 345 -45
rect 359 -47 361 -45
rect 386 -53 388 -36
rect 392 -39 394 -36
rect 408 -53 410 -36
rect 424 -39 426 -36
rect 50 -72 52 -70
rect 56 -72 58 -70
rect 72 -72 74 -70
rect 88 -72 90 -70
rect 94 -72 96 -70
rect 110 -72 112 -70
rect 131 -72 133 -70
rect 137 -72 139 -70
rect 153 -72 155 -70
rect 169 -72 171 -70
rect 175 -72 177 -70
rect 191 -72 193 -70
rect 218 -72 220 -55
rect 224 -58 226 -55
rect 240 -72 242 -55
rect 256 -58 258 -55
rect 218 -97 220 -76
rect 224 -97 226 -90
rect 240 -97 242 -76
rect 256 -97 258 -62
rect 262 -65 264 -55
rect 278 -72 280 -55
rect 299 -72 301 -55
rect 305 -58 307 -55
rect 321 -72 323 -55
rect 337 -58 339 -55
rect 262 -97 264 -83
rect 278 -97 280 -76
rect 299 -97 301 -76
rect 305 -97 307 -90
rect 321 -97 323 -76
rect 337 -97 339 -62
rect 343 -65 345 -55
rect 359 -72 361 -55
rect 343 -97 345 -83
rect 359 -97 361 -76
rect 386 -78 388 -57
rect 392 -78 394 -71
rect 408 -78 410 -57
rect 424 -78 426 -43
rect 430 -46 432 -36
rect 446 -53 448 -36
rect 467 -53 469 -36
rect 473 -39 475 -36
rect 489 -53 491 -36
rect 505 -39 507 -36
rect 430 -78 432 -64
rect 446 -78 448 -57
rect 467 -78 469 -57
rect 473 -78 475 -71
rect 489 -78 491 -57
rect 505 -78 507 -43
rect 511 -46 513 -36
rect 527 -53 529 -36
rect 511 -78 513 -64
rect 527 -78 529 -57
rect 386 -84 388 -82
rect 392 -84 394 -82
rect 408 -84 410 -82
rect 424 -84 426 -82
rect 430 -84 432 -82
rect 446 -84 448 -82
rect 467 -84 469 -82
rect 473 -84 475 -82
rect 489 -84 491 -82
rect 505 -84 507 -82
rect 511 -84 513 -82
rect 527 -84 529 -82
rect 218 -103 220 -101
rect 224 -103 226 -101
rect 240 -103 242 -101
rect 256 -103 258 -101
rect 262 -103 264 -101
rect 278 -103 280 -101
rect 299 -103 301 -101
rect 305 -103 307 -101
rect 321 -103 323 -101
rect 337 -103 339 -101
rect 343 -103 345 -101
rect 359 -103 361 -101
rect 445 -102 447 -98
rect 469 -102 471 -98
rect 445 -108 447 -106
rect 469 -108 471 -106
rect 465 -113 467 -111
rect 465 -120 467 -117
rect 218 -129 220 -127
rect 224 -129 226 -127
rect 240 -129 242 -127
rect 256 -129 258 -127
rect 262 -129 264 -127
rect 278 -129 280 -127
rect 299 -129 301 -127
rect 305 -129 307 -127
rect 321 -129 323 -127
rect 337 -129 339 -127
rect 343 -129 345 -127
rect 359 -129 361 -127
rect 453 -130 456 -129
rect 449 -131 456 -130
rect 460 -131 462 -129
rect 218 -154 220 -133
rect 224 -140 226 -133
rect 240 -154 242 -133
rect 218 -175 220 -158
rect 224 -175 226 -172
rect 240 -175 242 -158
rect 256 -168 258 -133
rect 262 -147 264 -133
rect 278 -154 280 -133
rect 299 -154 301 -133
rect 305 -140 307 -133
rect 321 -154 323 -133
rect 256 -175 258 -172
rect 262 -175 264 -165
rect 278 -175 280 -158
rect 299 -175 301 -158
rect 305 -175 307 -172
rect 321 -175 323 -158
rect 337 -168 339 -133
rect 343 -147 345 -133
rect 359 -154 361 -133
rect 445 -136 447 -134
rect 469 -136 471 -134
rect 445 -144 447 -140
rect 469 -144 471 -140
rect 337 -175 339 -172
rect 343 -175 345 -165
rect 359 -175 361 -158
rect 386 -160 388 -158
rect 392 -160 394 -158
rect 408 -160 410 -158
rect 424 -160 426 -158
rect 430 -160 432 -158
rect 446 -160 448 -158
rect 467 -160 469 -158
rect 473 -160 475 -158
rect 489 -160 491 -158
rect 505 -160 507 -158
rect 511 -160 513 -158
rect 527 -160 529 -158
rect 218 -185 220 -183
rect 224 -185 226 -183
rect 240 -185 242 -183
rect 256 -185 258 -183
rect 262 -185 264 -183
rect 278 -185 280 -183
rect 299 -185 301 -183
rect 305 -185 307 -183
rect 321 -185 323 -183
rect 337 -185 339 -183
rect 343 -185 345 -183
rect 359 -185 361 -183
rect 386 -185 388 -168
rect 392 -171 394 -168
rect 408 -185 410 -168
rect 424 -171 426 -168
rect 386 -210 388 -189
rect 392 -210 394 -203
rect 408 -210 410 -189
rect 424 -210 426 -175
rect 430 -178 432 -168
rect 446 -185 448 -168
rect 467 -185 469 -168
rect 473 -171 475 -168
rect 489 -185 491 -168
rect 505 -171 507 -168
rect 430 -210 432 -196
rect 446 -210 448 -189
rect 467 -210 469 -189
rect 473 -210 475 -203
rect 489 -210 491 -189
rect 505 -210 507 -175
rect 511 -178 513 -168
rect 527 -185 529 -168
rect 511 -210 513 -196
rect 527 -210 529 -189
rect 386 -216 388 -214
rect 392 -216 394 -214
rect 408 -216 410 -214
rect 424 -216 426 -214
rect 430 -216 432 -214
rect 446 -216 448 -214
rect 467 -216 469 -214
rect 473 -216 475 -214
rect 489 -216 491 -214
rect 505 -216 507 -214
rect 511 -216 513 -214
rect 527 -216 529 -214
rect 386 -226 388 -224
rect 392 -226 394 -224
rect 408 -226 410 -224
rect 424 -226 426 -224
rect 430 -226 432 -224
rect 446 -226 448 -224
rect 467 -226 469 -224
rect 473 -226 475 -224
rect 489 -226 491 -224
rect 505 -226 507 -224
rect 511 -226 513 -224
rect 527 -226 529 -224
rect 386 -251 388 -230
rect 392 -237 394 -230
rect 408 -251 410 -230
rect 386 -272 388 -255
rect 392 -272 394 -269
rect 408 -272 410 -255
rect 424 -265 426 -230
rect 430 -244 432 -230
rect 446 -251 448 -230
rect 467 -251 469 -230
rect 473 -237 475 -230
rect 489 -251 491 -230
rect 424 -272 426 -269
rect 430 -272 432 -262
rect 446 -272 448 -255
rect 467 -272 469 -255
rect 473 -272 475 -269
rect 489 -272 491 -255
rect 505 -265 507 -230
rect 511 -244 513 -230
rect 527 -251 529 -230
rect 505 -272 507 -269
rect 511 -272 513 -262
rect 527 -272 529 -255
rect 386 -282 388 -280
rect 392 -282 394 -280
rect 408 -282 410 -280
rect 424 -282 426 -280
rect 430 -282 432 -280
rect 446 -282 448 -280
rect 467 -282 469 -280
rect 473 -282 475 -280
rect 489 -282 491 -280
rect 505 -282 507 -280
rect 511 -282 513 -280
rect 527 -282 529 -280
<< polycontact >>
rect 55 183 59 187
rect 87 183 91 187
rect 49 169 53 173
rect 71 169 75 173
rect 55 155 59 159
rect 93 176 97 180
rect 136 183 140 187
rect 168 183 172 187
rect 109 169 113 173
rect 130 169 134 173
rect 152 169 156 173
rect 93 162 97 166
rect 136 155 140 159
rect 174 176 178 180
rect 190 169 194 173
rect 174 162 178 166
rect 108 128 112 132
rect 132 128 136 132
rect 128 102 132 106
rect 113 96 117 100
rect 108 78 112 82
rect 132 78 136 82
rect 223 70 227 74
rect 255 70 259 74
rect 55 51 59 55
rect 87 51 91 55
rect 49 37 53 41
rect 71 37 75 41
rect 55 23 59 27
rect 93 44 97 48
rect 136 51 140 55
rect 168 51 172 55
rect 109 37 113 41
rect 130 37 134 41
rect 152 37 156 41
rect 93 30 97 34
rect 136 23 140 27
rect 174 44 178 48
rect 217 56 221 60
rect 239 56 243 60
rect 190 37 194 41
rect 174 30 178 34
rect 223 42 227 46
rect 261 63 265 67
rect 304 70 308 74
rect 336 70 340 74
rect 277 56 281 60
rect 298 56 302 60
rect 320 56 324 60
rect 261 49 265 53
rect 304 42 308 46
rect 342 63 346 67
rect 358 56 362 60
rect 342 49 346 53
rect 276 15 280 19
rect 300 15 304 19
rect 296 -11 300 -7
rect 281 -17 285 -13
rect 55 -31 59 -27
rect 49 -45 53 -41
rect 71 -45 75 -41
rect 55 -59 59 -55
rect 93 -38 97 -34
rect 136 -31 140 -27
rect 109 -45 113 -41
rect 130 -45 134 -41
rect 152 -45 156 -41
rect 93 -52 97 -48
rect 87 -59 91 -55
rect 136 -59 140 -55
rect 174 -38 178 -34
rect 276 -35 280 -31
rect 300 -35 304 -31
rect 190 -45 194 -41
rect 174 -52 178 -48
rect 168 -59 172 -55
rect 391 -43 395 -39
rect 423 -43 427 -39
rect 223 -62 227 -58
rect 255 -62 259 -58
rect 217 -76 221 -72
rect 239 -76 243 -72
rect 223 -90 227 -86
rect 261 -69 265 -65
rect 304 -62 308 -58
rect 336 -62 340 -58
rect 277 -76 281 -72
rect 298 -76 302 -72
rect 320 -76 324 -72
rect 261 -83 265 -79
rect 304 -90 308 -86
rect 342 -69 346 -65
rect 385 -57 389 -53
rect 407 -57 411 -53
rect 358 -76 362 -72
rect 342 -83 346 -79
rect 391 -71 395 -67
rect 429 -50 433 -46
rect 472 -43 476 -39
rect 504 -43 508 -39
rect 445 -57 449 -53
rect 466 -57 470 -53
rect 488 -57 492 -53
rect 429 -64 433 -60
rect 472 -71 476 -67
rect 510 -50 514 -46
rect 526 -57 530 -53
rect 510 -64 514 -60
rect 444 -98 448 -94
rect 468 -98 472 -94
rect 464 -124 468 -120
rect 449 -130 453 -126
rect 223 -144 227 -140
rect 217 -158 221 -154
rect 239 -158 243 -154
rect 223 -172 227 -168
rect 261 -151 265 -147
rect 304 -144 308 -140
rect 277 -158 281 -154
rect 298 -158 302 -154
rect 320 -158 324 -154
rect 261 -165 265 -161
rect 255 -172 259 -168
rect 304 -172 308 -168
rect 342 -151 346 -147
rect 444 -148 448 -144
rect 468 -148 472 -144
rect 358 -158 362 -154
rect 342 -165 346 -161
rect 336 -172 340 -168
rect 391 -175 395 -171
rect 423 -175 427 -171
rect 385 -189 389 -185
rect 407 -189 411 -185
rect 391 -203 395 -199
rect 429 -182 433 -178
rect 472 -175 476 -171
rect 504 -175 508 -171
rect 445 -189 449 -185
rect 466 -189 470 -185
rect 488 -189 492 -185
rect 429 -196 433 -192
rect 472 -203 476 -199
rect 510 -182 514 -178
rect 526 -189 530 -185
rect 510 -196 514 -192
rect 391 -241 395 -237
rect 385 -255 389 -251
rect 407 -255 411 -251
rect 391 -269 395 -265
rect 429 -248 433 -244
rect 472 -241 476 -237
rect 445 -255 449 -251
rect 466 -255 470 -251
rect 488 -255 492 -251
rect 429 -262 433 -258
rect 423 -269 427 -265
rect 472 -269 476 -265
rect 510 -248 514 -244
rect 526 -255 530 -251
rect 510 -262 514 -258
rect 504 -269 508 -265
<< metal1 >>
rect 34 202 45 206
rect 49 202 61 206
rect 65 202 76 206
rect 80 202 98 206
rect 102 202 126 206
rect 130 202 142 206
rect 146 202 157 206
rect 161 202 179 206
rect 183 202 198 206
rect 45 198 49 202
rect 67 198 71 202
rect 83 198 87 202
rect 105 198 109 202
rect 126 198 130 202
rect 148 198 152 202
rect 164 198 168 202
rect 186 198 190 202
rect 45 183 55 187
rect 79 183 87 187
rect 131 183 136 187
rect 160 183 168 187
rect 38 176 93 180
rect 97 176 174 180
rect 45 169 49 173
rect 63 169 71 173
rect 75 169 97 173
rect 101 169 109 173
rect 125 169 130 173
rect 144 169 152 173
rect 156 169 178 173
rect 182 169 190 173
rect 45 162 93 166
rect 97 162 127 166
rect 131 162 174 166
rect 38 155 55 159
rect 59 155 136 159
rect 45 140 49 144
rect 67 140 71 144
rect 83 140 87 144
rect 105 140 109 144
rect 126 140 130 144
rect 148 140 152 144
rect 164 140 168 144
rect 186 140 190 144
rect 34 136 38 140
rect 42 136 80 140
rect 84 136 89 140
rect 93 136 101 140
rect 105 136 161 140
rect 165 136 170 140
rect 174 136 182 140
rect 186 136 198 140
rect 112 128 113 132
rect 136 128 194 132
rect 116 120 120 124
rect 124 120 128 124
rect 31 109 104 113
rect 108 109 124 113
rect 140 109 575 113
rect 132 102 186 106
rect 101 97 113 100
rect 116 86 120 90
rect 124 86 128 90
rect 202 89 213 93
rect 217 89 229 93
rect 233 89 244 93
rect 248 89 266 93
rect 270 89 294 93
rect 298 89 310 93
rect 314 89 325 93
rect 329 89 347 93
rect 351 89 366 93
rect 213 85 217 89
rect 235 85 239 89
rect 251 85 255 89
rect 273 85 277 89
rect 294 85 298 89
rect 316 85 320 89
rect 332 85 336 89
rect 354 85 358 89
rect 112 78 113 82
rect 136 78 194 82
rect 34 70 45 74
rect 49 70 61 74
rect 65 70 76 74
rect 80 70 126 74
rect 130 70 142 74
rect 146 70 157 74
rect 161 70 179 74
rect 183 70 198 74
rect 213 70 223 74
rect 247 70 255 74
rect 299 70 304 74
rect 328 70 336 74
rect 45 66 49 70
rect 67 66 71 70
rect 83 66 87 70
rect 105 66 109 70
rect 126 66 130 70
rect 148 66 152 70
rect 164 66 168 70
rect 186 66 190 70
rect 206 63 261 67
rect 265 63 342 67
rect 213 56 217 60
rect 231 56 239 60
rect 243 56 265 60
rect 269 56 277 60
rect 293 56 298 60
rect 312 56 320 60
rect 324 56 346 60
rect 350 56 358 60
rect 45 51 55 55
rect 79 51 87 55
rect 131 51 136 55
rect 160 51 168 55
rect 213 49 261 53
rect 265 49 295 53
rect 299 49 342 53
rect 38 44 93 48
rect 97 44 174 48
rect 206 42 223 46
rect 227 42 304 46
rect 45 37 49 41
rect 63 37 71 41
rect 75 37 97 41
rect 101 37 109 41
rect 125 37 130 41
rect 144 37 152 41
rect 156 37 178 41
rect 182 37 190 41
rect 45 30 93 34
rect 97 30 127 34
rect 131 30 174 34
rect 213 27 217 31
rect 235 27 239 31
rect 251 27 255 31
rect 273 27 277 31
rect 294 27 298 31
rect 316 27 320 31
rect 332 27 336 31
rect 354 27 358 31
rect 38 23 55 27
rect 59 23 136 27
rect 202 23 206 27
rect 210 23 248 27
rect 252 23 257 27
rect 261 23 269 27
rect 273 23 329 27
rect 333 23 338 27
rect 342 23 350 27
rect 354 23 366 27
rect 280 15 281 19
rect 304 15 362 19
rect 45 8 49 12
rect 67 8 71 12
rect 83 8 87 12
rect 105 8 109 12
rect 126 8 130 12
rect 148 8 152 12
rect 164 8 168 12
rect 186 8 190 12
rect 34 4 112 8
rect 116 4 143 8
rect 147 4 195 8
rect 284 7 288 11
rect 292 7 296 11
rect 31 -4 272 0
rect 276 -4 292 0
rect 308 -4 580 0
rect 34 -12 38 -8
rect 42 -12 80 -8
rect 84 -12 89 -8
rect 93 -12 101 -8
rect 105 -12 161 -8
rect 165 -12 170 -8
rect 174 -12 182 -8
rect 186 -12 198 -8
rect 300 -11 354 -7
rect 45 -16 49 -12
rect 67 -16 71 -12
rect 83 -16 87 -12
rect 105 -16 109 -12
rect 126 -16 130 -12
rect 148 -16 152 -12
rect 164 -16 168 -12
rect 186 -16 190 -12
rect 269 -16 281 -13
rect 284 -27 288 -23
rect 292 -27 296 -23
rect 370 -24 381 -20
rect 385 -24 397 -20
rect 401 -24 412 -20
rect 416 -24 434 -20
rect 438 -24 462 -20
rect 466 -24 478 -20
rect 482 -24 493 -20
rect 497 -24 515 -20
rect 519 -24 534 -20
rect 38 -31 55 -27
rect 59 -31 136 -27
rect 381 -28 385 -24
rect 403 -28 407 -24
rect 419 -28 423 -24
rect 441 -28 445 -24
rect 462 -28 466 -24
rect 484 -28 488 -24
rect 500 -28 504 -24
rect 522 -28 526 -24
rect 45 -38 93 -34
rect 97 -38 127 -34
rect 131 -38 174 -34
rect 280 -35 281 -31
rect 304 -35 362 -31
rect 45 -45 49 -41
rect 63 -45 71 -41
rect 75 -45 97 -41
rect 101 -45 109 -41
rect 125 -45 130 -41
rect 144 -45 152 -41
rect 156 -45 178 -41
rect 182 -45 190 -41
rect 202 -43 213 -39
rect 217 -43 229 -39
rect 233 -43 244 -39
rect 248 -43 294 -39
rect 298 -43 310 -39
rect 314 -43 325 -39
rect 329 -43 347 -39
rect 351 -43 366 -39
rect 381 -43 391 -39
rect 415 -43 423 -39
rect 467 -43 472 -39
rect 496 -43 504 -39
rect 213 -47 217 -43
rect 235 -47 239 -43
rect 251 -47 255 -43
rect 273 -47 277 -43
rect 294 -47 298 -43
rect 316 -47 320 -43
rect 332 -47 336 -43
rect 354 -47 358 -43
rect 38 -52 93 -48
rect 97 -52 174 -48
rect 374 -50 429 -46
rect 433 -50 510 -46
rect 45 -59 55 -55
rect 79 -59 87 -55
rect 131 -59 136 -55
rect 160 -59 168 -55
rect 381 -57 385 -53
rect 399 -57 407 -53
rect 411 -57 433 -53
rect 437 -57 445 -53
rect 461 -57 466 -53
rect 480 -57 488 -53
rect 492 -57 514 -53
rect 518 -57 526 -53
rect 213 -62 223 -58
rect 247 -62 255 -58
rect 299 -62 304 -58
rect 328 -62 336 -58
rect 381 -64 429 -60
rect 433 -64 463 -60
rect 467 -64 510 -60
rect 206 -69 261 -65
rect 265 -69 342 -65
rect 45 -74 49 -70
rect 67 -74 71 -70
rect 83 -74 87 -70
rect 105 -74 109 -70
rect 126 -74 130 -70
rect 148 -74 152 -70
rect 164 -74 168 -70
rect 186 -74 190 -70
rect 374 -71 391 -67
rect 395 -71 472 -67
rect 34 -78 45 -74
rect 49 -78 61 -74
rect 65 -78 76 -74
rect 80 -78 126 -74
rect 130 -78 142 -74
rect 146 -78 157 -74
rect 161 -78 179 -74
rect 183 -78 198 -74
rect 213 -76 217 -72
rect 231 -76 239 -72
rect 243 -76 265 -72
rect 269 -76 277 -72
rect 293 -76 298 -72
rect 312 -76 320 -72
rect 324 -76 346 -72
rect 350 -76 358 -72
rect 213 -83 261 -79
rect 265 -83 295 -79
rect 299 -83 342 -79
rect 381 -86 385 -82
rect 403 -86 407 -82
rect 419 -86 423 -82
rect 441 -86 445 -82
rect 462 -86 466 -82
rect 484 -86 488 -82
rect 500 -86 504 -82
rect 522 -86 526 -82
rect 206 -90 223 -86
rect 227 -90 304 -86
rect 370 -90 374 -86
rect 378 -90 416 -86
rect 420 -90 425 -86
rect 429 -90 437 -86
rect 441 -90 497 -86
rect 501 -90 506 -86
rect 510 -90 518 -86
rect 522 -90 534 -86
rect 448 -98 449 -94
rect 472 -98 530 -94
rect 213 -105 217 -101
rect 235 -105 239 -101
rect 251 -105 255 -101
rect 273 -105 277 -101
rect 294 -105 298 -101
rect 316 -105 320 -101
rect 332 -105 336 -101
rect 354 -105 358 -101
rect 202 -109 280 -105
rect 284 -109 311 -105
rect 315 -109 363 -105
rect 452 -106 456 -102
rect 460 -106 464 -102
rect 30 -117 440 -113
rect 444 -117 460 -113
rect 476 -117 596 -113
rect 202 -125 206 -121
rect 210 -125 248 -121
rect 252 -125 257 -121
rect 261 -125 269 -121
rect 273 -125 329 -121
rect 333 -125 338 -121
rect 342 -125 350 -121
rect 354 -125 366 -121
rect 468 -124 522 -120
rect 213 -129 217 -125
rect 235 -129 239 -125
rect 251 -129 255 -125
rect 273 -129 277 -125
rect 294 -129 298 -125
rect 316 -129 320 -125
rect 332 -129 336 -125
rect 354 -129 358 -125
rect 437 -129 449 -126
rect 452 -140 456 -136
rect 460 -140 464 -136
rect 206 -144 223 -140
rect 227 -144 304 -140
rect 213 -151 261 -147
rect 265 -151 295 -147
rect 299 -151 342 -147
rect 448 -148 449 -144
rect 472 -148 530 -144
rect 213 -158 217 -154
rect 231 -158 239 -154
rect 243 -158 265 -154
rect 269 -158 277 -154
rect 293 -158 298 -154
rect 312 -158 320 -154
rect 324 -158 346 -154
rect 350 -158 358 -154
rect 370 -156 381 -152
rect 385 -156 397 -152
rect 401 -156 412 -152
rect 416 -156 462 -152
rect 466 -156 478 -152
rect 482 -156 493 -152
rect 497 -156 515 -152
rect 519 -156 534 -152
rect 381 -160 385 -156
rect 403 -160 407 -156
rect 419 -160 423 -156
rect 441 -160 445 -156
rect 462 -160 466 -156
rect 484 -160 488 -156
rect 500 -160 504 -156
rect 522 -160 526 -156
rect 206 -165 261 -161
rect 265 -165 342 -161
rect 213 -172 223 -168
rect 247 -172 255 -168
rect 299 -172 304 -168
rect 328 -172 336 -168
rect 381 -175 391 -171
rect 415 -175 423 -171
rect 467 -175 472 -171
rect 496 -175 504 -171
rect 374 -182 429 -178
rect 433 -182 510 -178
rect 213 -187 217 -183
rect 235 -187 239 -183
rect 251 -187 255 -183
rect 273 -187 277 -183
rect 294 -187 298 -183
rect 316 -187 320 -183
rect 332 -187 336 -183
rect 354 -187 358 -183
rect 202 -191 213 -187
rect 217 -191 229 -187
rect 233 -191 244 -187
rect 248 -191 294 -187
rect 298 -191 310 -187
rect 314 -191 325 -187
rect 329 -191 347 -187
rect 351 -191 366 -187
rect 381 -189 385 -185
rect 399 -189 407 -185
rect 411 -189 433 -185
rect 437 -189 445 -185
rect 461 -189 466 -185
rect 480 -189 488 -185
rect 492 -189 514 -185
rect 518 -189 526 -185
rect 381 -196 429 -192
rect 433 -196 463 -192
rect 467 -196 510 -192
rect 374 -203 391 -199
rect 395 -203 472 -199
rect 381 -218 385 -214
rect 403 -218 407 -214
rect 419 -218 423 -214
rect 441 -218 445 -214
rect 462 -218 466 -214
rect 484 -218 488 -214
rect 500 -218 504 -214
rect 522 -218 526 -214
rect 370 -222 374 -218
rect 378 -222 416 -218
rect 420 -222 425 -218
rect 429 -222 437 -218
rect 441 -222 448 -218
rect 452 -222 479 -218
rect 483 -222 497 -218
rect 501 -222 506 -218
rect 510 -222 518 -218
rect 522 -222 534 -218
rect 381 -226 385 -222
rect 403 -226 407 -222
rect 419 -226 423 -222
rect 441 -226 445 -222
rect 462 -226 466 -222
rect 484 -226 488 -222
rect 500 -226 504 -222
rect 522 -226 526 -222
rect 374 -241 391 -237
rect 395 -241 472 -237
rect 381 -248 429 -244
rect 433 -248 463 -244
rect 467 -248 510 -244
rect 381 -255 385 -251
rect 399 -255 407 -251
rect 411 -255 433 -251
rect 437 -255 445 -251
rect 461 -255 466 -251
rect 480 -255 488 -251
rect 492 -255 514 -251
rect 518 -255 526 -251
rect 374 -262 429 -258
rect 433 -262 510 -258
rect 381 -269 391 -265
rect 415 -269 423 -265
rect 467 -269 472 -265
rect 496 -269 504 -265
rect 381 -284 385 -280
rect 403 -284 407 -280
rect 419 -284 423 -280
rect 441 -284 445 -280
rect 462 -284 466 -280
rect 484 -284 488 -280
rect 500 -284 504 -280
rect 522 -284 526 -280
rect 370 -288 381 -284
rect 385 -288 397 -284
rect 401 -288 412 -284
rect 416 -288 462 -284
rect 466 -288 478 -284
rect 482 -288 493 -284
rect 497 -288 515 -284
rect 519 -288 534 -284
<< m2contact >>
rect 59 190 63 194
rect 75 190 79 194
rect 97 190 101 194
rect 113 190 117 194
rect 140 190 144 194
rect 156 190 160 194
rect 178 190 182 194
rect 194 190 198 194
rect 41 183 45 187
rect 75 183 79 187
rect 127 183 131 187
rect 156 183 160 187
rect 34 176 38 180
rect 59 169 63 173
rect 97 169 101 173
rect 140 169 144 173
rect 178 169 182 173
rect 41 162 45 166
rect 127 162 131 166
rect 34 155 38 159
rect 59 148 63 152
rect 75 148 79 152
rect 97 148 101 152
rect 113 148 117 152
rect 140 148 144 152
rect 156 148 160 152
rect 178 148 182 152
rect 194 148 198 152
rect 113 128 117 132
rect 194 128 198 132
rect 120 120 124 124
rect 104 116 108 120
rect 136 116 140 120
rect 104 109 108 113
rect 136 109 140 113
rect 120 102 124 106
rect 186 102 190 106
rect 97 96 101 100
rect 104 90 108 94
rect 136 90 140 94
rect 120 86 124 90
rect 113 78 117 82
rect 194 78 198 82
rect 227 77 231 81
rect 243 77 247 81
rect 265 77 269 81
rect 281 77 285 81
rect 308 77 312 81
rect 324 77 328 81
rect 346 77 350 81
rect 362 77 366 81
rect 209 70 213 74
rect 243 70 247 74
rect 295 70 299 74
rect 324 70 328 74
rect 59 58 63 62
rect 75 58 79 62
rect 97 58 101 62
rect 113 58 117 62
rect 140 58 144 62
rect 156 58 160 62
rect 178 58 182 62
rect 202 63 206 67
rect 194 58 198 62
rect 227 56 231 60
rect 265 56 269 60
rect 308 56 312 60
rect 346 56 350 60
rect 41 51 45 55
rect 75 51 79 55
rect 127 51 131 55
rect 156 51 160 55
rect 209 49 213 53
rect 295 49 299 53
rect 34 44 38 48
rect 202 42 206 46
rect 59 37 63 41
rect 97 37 101 41
rect 140 37 144 41
rect 178 37 182 41
rect 227 35 231 39
rect 243 35 247 39
rect 265 35 269 39
rect 281 35 285 39
rect 308 35 312 39
rect 324 35 328 39
rect 346 35 350 39
rect 362 35 366 39
rect 41 30 45 34
rect 127 30 131 34
rect 34 23 38 27
rect 59 16 63 20
rect 75 16 79 20
rect 97 16 101 20
rect 113 16 117 20
rect 140 16 144 20
rect 156 16 160 20
rect 178 16 182 20
rect 194 16 198 20
rect 281 15 285 19
rect 362 15 366 19
rect 288 7 292 11
rect 272 3 276 7
rect 304 3 308 7
rect 272 -4 276 0
rect 304 -4 308 0
rect 288 -11 292 -7
rect 354 -11 358 -7
rect 265 -17 269 -13
rect 59 -24 63 -20
rect 75 -24 79 -20
rect 97 -24 101 -20
rect 113 -24 117 -20
rect 140 -24 144 -20
rect 156 -24 160 -20
rect 178 -24 182 -20
rect 194 -24 198 -20
rect 272 -23 276 -19
rect 304 -23 308 -19
rect 288 -27 292 -23
rect 34 -31 38 -27
rect 41 -38 45 -34
rect 127 -38 131 -34
rect 281 -35 285 -31
rect 362 -35 366 -31
rect 395 -36 399 -32
rect 411 -36 415 -32
rect 433 -36 437 -32
rect 449 -36 453 -32
rect 476 -36 480 -32
rect 492 -36 496 -32
rect 514 -36 518 -32
rect 530 -36 534 -32
rect 59 -45 63 -41
rect 97 -45 101 -41
rect 140 -45 144 -41
rect 178 -45 182 -41
rect 377 -43 381 -39
rect 411 -43 415 -39
rect 463 -43 467 -39
rect 492 -43 496 -39
rect 34 -52 38 -48
rect 227 -55 231 -51
rect 243 -55 247 -51
rect 265 -55 269 -51
rect 281 -55 285 -51
rect 308 -55 312 -51
rect 324 -55 328 -51
rect 346 -55 350 -51
rect 370 -50 374 -46
rect 362 -55 366 -51
rect 41 -59 45 -55
rect 75 -59 79 -55
rect 127 -59 131 -55
rect 156 -59 160 -55
rect 395 -57 399 -53
rect 433 -57 437 -53
rect 476 -57 480 -53
rect 514 -57 518 -53
rect 209 -62 213 -58
rect 243 -62 247 -58
rect 295 -62 299 -58
rect 324 -62 328 -58
rect 59 -66 63 -62
rect 75 -66 79 -62
rect 97 -66 101 -62
rect 113 -66 117 -62
rect 140 -66 144 -62
rect 156 -66 160 -62
rect 178 -66 182 -62
rect 194 -66 198 -62
rect 377 -64 381 -60
rect 463 -64 467 -60
rect 202 -69 206 -65
rect 370 -71 374 -67
rect 227 -76 231 -72
rect 265 -76 269 -72
rect 308 -76 312 -72
rect 346 -76 350 -72
rect 395 -78 399 -74
rect 411 -78 415 -74
rect 433 -78 437 -74
rect 449 -78 453 -74
rect 476 -78 480 -74
rect 492 -78 496 -74
rect 514 -78 518 -74
rect 530 -78 534 -74
rect 209 -83 213 -79
rect 295 -83 299 -79
rect 202 -90 206 -86
rect 227 -97 231 -93
rect 243 -97 247 -93
rect 265 -97 269 -93
rect 281 -97 285 -93
rect 308 -97 312 -93
rect 324 -97 328 -93
rect 346 -97 350 -93
rect 362 -97 366 -93
rect 449 -98 453 -94
rect 530 -98 534 -94
rect 456 -106 460 -102
rect 440 -110 444 -106
rect 472 -110 476 -106
rect 440 -117 444 -113
rect 472 -117 476 -113
rect 456 -124 460 -120
rect 522 -124 526 -120
rect 433 -130 437 -126
rect 227 -137 231 -133
rect 243 -137 247 -133
rect 265 -137 269 -133
rect 281 -137 285 -133
rect 308 -137 312 -133
rect 324 -137 328 -133
rect 346 -137 350 -133
rect 362 -137 366 -133
rect 440 -136 444 -132
rect 472 -136 476 -132
rect 456 -140 460 -136
rect 202 -144 206 -140
rect 209 -151 213 -147
rect 295 -151 299 -147
rect 449 -148 453 -144
rect 530 -148 534 -144
rect 227 -158 231 -154
rect 265 -158 269 -154
rect 308 -158 312 -154
rect 346 -158 350 -154
rect 202 -165 206 -161
rect 395 -168 399 -164
rect 411 -168 415 -164
rect 433 -168 437 -164
rect 449 -168 453 -164
rect 476 -168 480 -164
rect 492 -168 496 -164
rect 514 -168 518 -164
rect 530 -168 534 -164
rect 209 -172 213 -168
rect 243 -172 247 -168
rect 295 -172 299 -168
rect 324 -172 328 -168
rect 377 -175 381 -171
rect 411 -175 415 -171
rect 463 -175 467 -171
rect 492 -175 496 -171
rect 227 -179 231 -175
rect 243 -179 247 -175
rect 265 -179 269 -175
rect 281 -179 285 -175
rect 308 -179 312 -175
rect 324 -179 328 -175
rect 346 -179 350 -175
rect 362 -179 366 -175
rect 370 -182 374 -178
rect 395 -189 399 -185
rect 433 -189 437 -185
rect 476 -189 480 -185
rect 514 -189 518 -185
rect 377 -196 381 -192
rect 463 -196 467 -192
rect 370 -203 374 -199
rect 395 -210 399 -206
rect 411 -210 415 -206
rect 433 -210 437 -206
rect 449 -210 453 -206
rect 476 -210 480 -206
rect 492 -210 496 -206
rect 514 -210 518 -206
rect 530 -210 534 -206
rect 395 -234 399 -230
rect 411 -234 415 -230
rect 433 -234 437 -230
rect 449 -234 453 -230
rect 476 -234 480 -230
rect 492 -234 496 -230
rect 514 -234 518 -230
rect 530 -234 534 -230
rect 370 -241 374 -237
rect 377 -248 381 -244
rect 463 -248 467 -244
rect 395 -255 399 -251
rect 433 -255 437 -251
rect 476 -255 480 -251
rect 514 -255 518 -251
rect 370 -262 374 -258
rect 377 -269 381 -265
rect 411 -269 415 -265
rect 463 -269 467 -265
rect 492 -269 496 -265
rect 395 -276 399 -272
rect 411 -276 415 -272
rect 433 -276 437 -272
rect 449 -276 453 -272
rect 476 -276 480 -272
rect 492 -276 496 -272
rect 514 -276 518 -272
rect 530 -276 534 -272
<< metal2 >>
rect 34 180 38 206
rect 34 159 38 176
rect 34 48 38 155
rect 34 27 38 44
rect 34 -27 38 23
rect 34 -48 38 -31
rect 34 -78 38 -52
rect 41 187 45 206
rect 41 166 45 183
rect 41 55 45 162
rect 59 194 63 198
rect 59 173 63 190
rect 59 152 63 169
rect 59 144 63 148
rect 75 194 79 198
rect 75 187 79 190
rect 75 152 79 183
rect 75 144 79 148
rect 97 194 101 198
rect 97 173 101 190
rect 97 152 101 169
rect 97 144 101 148
rect 113 194 117 198
rect 113 152 117 190
rect 113 132 117 148
rect 120 124 124 212
rect 140 194 144 198
rect 127 166 131 183
rect 140 173 144 190
rect 140 152 144 169
rect 140 144 144 148
rect 156 194 160 198
rect 156 187 160 190
rect 156 152 160 183
rect 156 144 160 148
rect 178 194 182 198
rect 178 173 182 190
rect 178 152 182 169
rect 178 144 182 148
rect 194 194 198 198
rect 194 152 198 190
rect 194 132 198 148
rect 104 113 108 116
rect 97 74 101 96
rect 104 94 108 109
rect 120 106 124 120
rect 136 120 140 124
rect 136 113 140 116
rect 136 94 140 109
rect 136 86 140 90
rect 97 70 109 74
rect 41 34 45 51
rect 41 -34 45 30
rect 59 62 63 66
rect 59 41 63 58
rect 59 20 63 37
rect 59 12 63 16
rect 75 62 79 66
rect 75 55 79 58
rect 75 20 79 51
rect 75 12 79 16
rect 97 62 101 66
rect 97 41 101 58
rect 97 20 101 37
rect 97 12 101 16
rect 105 -8 109 70
rect 113 62 117 78
rect 113 20 117 58
rect 113 12 117 16
rect 105 -12 117 -8
rect 41 -55 45 -38
rect 41 -78 45 -59
rect 59 -20 63 -16
rect 59 -41 63 -24
rect 59 -62 63 -45
rect 59 -70 63 -66
rect 75 -20 79 -16
rect 75 -55 79 -24
rect 75 -62 79 -59
rect 75 -70 79 -66
rect 97 -20 101 -16
rect 97 -41 101 -24
rect 97 -62 101 -45
rect 97 -70 101 -66
rect 113 -20 117 -12
rect 113 -62 117 -24
rect 113 -70 117 -66
rect 120 -323 124 86
rect 140 62 144 66
rect 127 34 131 51
rect 140 41 144 58
rect 140 20 144 37
rect 140 12 144 16
rect 156 62 160 66
rect 156 55 160 58
rect 156 20 160 51
rect 156 12 160 16
rect 178 62 182 66
rect 178 41 182 58
rect 178 20 182 37
rect 178 12 182 16
rect 186 -8 190 102
rect 194 62 198 78
rect 194 20 198 58
rect 194 12 198 16
rect 202 67 206 93
rect 202 46 206 63
rect 186 -12 198 -8
rect 140 -20 144 -16
rect 127 -55 131 -38
rect 140 -41 144 -24
rect 140 -62 144 -45
rect 140 -70 144 -66
rect 156 -20 160 -16
rect 156 -55 160 -24
rect 156 -62 160 -59
rect 156 -70 160 -66
rect 178 -20 182 -16
rect 178 -41 182 -24
rect 178 -62 182 -45
rect 178 -70 182 -66
rect 194 -20 198 -12
rect 194 -62 198 -24
rect 194 -78 198 -66
rect 202 -65 206 42
rect 202 -86 206 -69
rect 202 -140 206 -90
rect 202 -161 206 -144
rect 202 -191 206 -165
rect 209 74 213 93
rect 209 53 213 70
rect 209 -58 213 49
rect 227 81 231 85
rect 227 60 231 77
rect 227 39 231 56
rect 227 31 231 35
rect 243 81 247 85
rect 243 74 247 77
rect 243 39 247 70
rect 243 31 247 35
rect 265 81 269 85
rect 265 60 269 77
rect 265 39 269 56
rect 265 31 269 35
rect 281 81 285 85
rect 281 39 285 77
rect 281 19 285 35
rect 288 11 292 243
rect 308 81 312 85
rect 295 53 299 70
rect 308 60 312 77
rect 308 39 312 56
rect 308 31 312 35
rect 324 81 328 85
rect 324 74 328 77
rect 324 39 328 70
rect 324 31 328 35
rect 346 81 350 85
rect 346 60 350 77
rect 346 39 350 56
rect 346 31 350 35
rect 362 81 366 85
rect 362 39 366 77
rect 362 19 366 35
rect 272 0 276 3
rect 265 -39 269 -17
rect 272 -19 276 -4
rect 288 -7 292 7
rect 304 7 308 11
rect 304 0 308 3
rect 304 -19 308 -4
rect 304 -27 308 -23
rect 265 -43 277 -39
rect 209 -79 213 -62
rect 209 -147 213 -83
rect 227 -51 231 -47
rect 227 -72 231 -55
rect 227 -93 231 -76
rect 227 -101 231 -97
rect 243 -51 247 -47
rect 243 -58 247 -55
rect 243 -93 247 -62
rect 243 -101 247 -97
rect 265 -51 269 -47
rect 265 -72 269 -55
rect 265 -93 269 -76
rect 265 -101 269 -97
rect 273 -121 277 -43
rect 281 -51 285 -35
rect 281 -93 285 -55
rect 281 -101 285 -97
rect 273 -125 285 -121
rect 209 -168 213 -151
rect 209 -191 213 -172
rect 227 -133 231 -129
rect 227 -154 231 -137
rect 227 -175 231 -158
rect 227 -183 231 -179
rect 243 -133 247 -129
rect 243 -168 247 -137
rect 243 -175 247 -172
rect 243 -183 247 -179
rect 265 -133 269 -129
rect 265 -154 269 -137
rect 265 -175 269 -158
rect 265 -183 269 -179
rect 281 -133 285 -125
rect 281 -175 285 -137
rect 281 -183 285 -179
rect 288 -314 292 -27
rect 308 -51 312 -47
rect 295 -79 299 -62
rect 308 -72 312 -55
rect 308 -93 312 -76
rect 308 -101 312 -97
rect 324 -51 328 -47
rect 324 -58 328 -55
rect 324 -93 328 -62
rect 324 -101 328 -97
rect 346 -51 350 -47
rect 346 -72 350 -55
rect 346 -93 350 -76
rect 346 -101 350 -97
rect 354 -121 358 -11
rect 362 -51 366 -35
rect 362 -93 366 -55
rect 362 -101 366 -97
rect 370 -46 374 -20
rect 370 -67 374 -50
rect 354 -125 366 -121
rect 308 -133 312 -129
rect 295 -168 299 -151
rect 308 -154 312 -137
rect 308 -175 312 -158
rect 308 -183 312 -179
rect 324 -133 328 -129
rect 324 -168 328 -137
rect 324 -175 328 -172
rect 324 -183 328 -179
rect 346 -133 350 -129
rect 346 -154 350 -137
rect 346 -175 350 -158
rect 346 -183 350 -179
rect 362 -133 366 -125
rect 362 -175 366 -137
rect 362 -191 366 -179
rect 370 -178 374 -71
rect 370 -199 374 -182
rect 370 -237 374 -203
rect 370 -258 374 -241
rect 370 -288 374 -262
rect 377 -39 381 -20
rect 377 -60 381 -43
rect 377 -171 381 -64
rect 395 -32 399 -28
rect 395 -53 399 -36
rect 395 -74 399 -57
rect 395 -82 399 -78
rect 411 -32 415 -28
rect 411 -39 415 -36
rect 411 -74 415 -43
rect 411 -82 415 -78
rect 433 -32 437 -28
rect 433 -53 437 -36
rect 433 -74 437 -57
rect 433 -82 437 -78
rect 449 -32 453 -28
rect 449 -74 453 -36
rect 449 -94 453 -78
rect 456 -102 460 227
rect 476 -32 480 -28
rect 463 -60 467 -43
rect 476 -53 480 -36
rect 476 -74 480 -57
rect 476 -82 480 -78
rect 492 -32 496 -28
rect 492 -39 496 -36
rect 492 -74 496 -43
rect 492 -82 496 -78
rect 514 -32 518 -28
rect 514 -53 518 -36
rect 514 -74 518 -57
rect 514 -82 518 -78
rect 530 -32 534 -28
rect 530 -74 534 -36
rect 530 -94 534 -78
rect 440 -113 444 -110
rect 433 -152 437 -130
rect 440 -132 444 -117
rect 456 -120 460 -106
rect 472 -106 476 -102
rect 472 -113 476 -110
rect 472 -132 476 -117
rect 472 -140 476 -136
rect 433 -156 445 -152
rect 377 -192 381 -175
rect 377 -244 381 -196
rect 395 -164 399 -160
rect 395 -185 399 -168
rect 395 -206 399 -189
rect 395 -214 399 -210
rect 411 -164 415 -160
rect 411 -171 415 -168
rect 411 -206 415 -175
rect 411 -214 415 -210
rect 433 -164 437 -160
rect 433 -185 437 -168
rect 433 -206 437 -189
rect 433 -214 437 -210
rect 441 -218 445 -156
rect 449 -164 453 -148
rect 449 -206 453 -168
rect 449 -214 453 -210
rect 441 -222 453 -218
rect 377 -265 381 -248
rect 377 -288 381 -269
rect 395 -230 399 -226
rect 395 -251 399 -234
rect 395 -272 399 -255
rect 395 -280 399 -276
rect 411 -230 415 -226
rect 411 -265 415 -234
rect 411 -272 415 -269
rect 411 -280 415 -276
rect 433 -230 437 -226
rect 433 -251 437 -234
rect 433 -272 437 -255
rect 433 -280 437 -276
rect 449 -230 453 -222
rect 449 -272 453 -234
rect 449 -280 453 -276
rect 456 -311 460 -140
rect 476 -164 480 -160
rect 463 -192 467 -175
rect 476 -185 480 -168
rect 476 -206 480 -189
rect 476 -214 480 -210
rect 492 -164 496 -160
rect 492 -171 496 -168
rect 492 -206 496 -175
rect 492 -214 496 -210
rect 514 -164 518 -160
rect 514 -185 518 -168
rect 514 -206 518 -189
rect 514 -214 518 -210
rect 522 -218 526 -124
rect 530 -164 534 -148
rect 530 -206 534 -168
rect 530 -214 534 -210
rect 522 -222 534 -218
rect 476 -230 480 -226
rect 463 -265 467 -248
rect 476 -251 480 -234
rect 476 -272 480 -255
rect 476 -280 480 -276
rect 492 -230 496 -226
rect 492 -265 496 -234
rect 492 -272 496 -269
rect 492 -280 496 -276
rect 514 -230 518 -226
rect 514 -251 518 -234
rect 514 -272 518 -255
rect 514 -280 518 -276
rect 530 -230 534 -222
rect 530 -272 534 -234
rect 530 -288 534 -276
<< labels >>
rlabel metal1 46 -44 46 -44 1 in5
rlabel metal1 126 -43 126 -43 1 in6
rlabel metal2 115 -44 115 -44 1 out5
rlabel metal2 196 -43 196 -43 1 out6
rlabel metal1 134 -10 134 -10 5 GND!
rlabel metal1 136 -76 136 -76 5 Vdd!
rlabel metal1 53 -10 53 -10 5 GND!
rlabel metal1 55 -76 55 -76 5 Vdd!
rlabel metal1 192 6 192 6 1 GND!
rlabel polysilicon 119 96 119 96 1 5
rlabel polysilicon 130 108 130 108 1 6
rlabel polysilicon 134 84 134 84 1 4
rlabel metal2 196 39 196 39 1 out4
rlabel metal1 126 39 126 39 1 in4
rlabel metal1 136 72 136 72 1 Vdd!
rlabel polysilicon 110 84 110 84 1 3
rlabel metal2 115 39 115 39 1 out3
rlabel metal1 47 39 47 39 1 in3
rlabel metal1 55 72 55 72 1 Vdd!
rlabel polysilicon 110 126 110 126 1 1
rlabel polysilicon 134 126 134 126 1 2
rlabel metal2 196 171 196 171 1 out2
rlabel metal1 126 170 126 170 1 in2
rlabel metal1 134 138 134 138 1 GND!
rlabel metal1 136 204 136 204 1 Vdd!
rlabel metal2 43 171 43 171 1 clk_b
rlabel metal2 37 169 37 169 3 clk
rlabel metal2 115 171 115 171 1 out1
rlabel metal1 53 138 53 138 1 GND!
rlabel metal1 47 171 47 171 1 in1
rlabel metal1 55 204 55 204 1 Vdd!
rlabel metal1 97 111 97 111 1 A
rlabel metal2 122 131 122 131 1 B
rlabel metal1 155 111 155 111 1 C
rlabel metal2 122 79 122 79 1 D
<< end >>
