magic
tech scmos
timestamp 1608229708
<< ntransistor >>
rect 8 564 10 568
rect 13 564 15 568
rect 29 564 31 568
rect 45 564 47 568
rect 50 564 52 568
rect 71 564 73 568
rect 87 564 89 568
rect 103 564 105 568
rect 108 564 110 568
rect 124 564 126 568
rect 140 564 142 568
rect 145 564 147 568
rect 161 564 163 568
rect 177 564 179 568
rect 182 564 184 568
rect 203 564 205 568
rect 219 564 221 568
rect 235 564 237 568
rect 240 564 242 568
rect 256 564 258 568
rect 272 564 274 568
rect 277 564 279 568
rect 293 564 295 568
rect 309 564 311 568
rect 314 564 316 568
rect 335 564 337 568
rect 351 564 353 568
rect 367 564 369 568
rect 372 564 374 568
rect 388 564 390 568
rect 404 564 406 568
rect 409 564 411 568
rect 425 564 427 568
rect 441 564 443 568
rect 446 564 448 568
rect 467 564 469 568
rect 483 564 485 568
rect 499 564 501 568
rect 504 564 506 568
rect 520 564 522 568
rect 187 498 189 502
rect 213 494 215 498
rect 218 494 220 498
rect 268 498 270 502
rect 294 494 296 498
rect 299 494 301 498
rect 241 490 243 494
rect 13 485 15 489
rect 29 485 31 489
rect 45 485 47 489
rect 68 485 70 489
rect 73 485 75 489
rect 99 485 101 489
rect 120 485 122 489
rect 140 485 142 489
rect 145 485 147 489
rect 163 485 165 489
rect 322 490 324 494
rect 13 439 15 443
rect 29 439 31 443
rect 45 439 47 443
rect 68 439 70 443
rect 73 439 75 443
rect 99 439 101 443
rect 120 439 122 443
rect 140 439 142 443
rect 145 439 147 443
rect 163 439 165 443
rect 213 438 215 442
rect 218 438 220 442
rect 294 438 296 442
rect 299 438 301 442
rect 213 362 215 366
rect 218 362 220 366
rect 292 366 294 370
rect 318 362 320 366
rect 323 362 325 366
rect 241 358 243 362
rect 13 353 15 357
rect 29 353 31 357
rect 45 353 47 357
rect 68 353 70 357
rect 73 353 75 357
rect 99 353 101 357
rect 120 353 122 357
rect 140 353 142 357
rect 145 353 147 357
rect 163 353 165 357
rect 346 358 348 362
rect 13 307 15 311
rect 29 307 31 311
rect 45 307 47 311
rect 68 307 70 311
rect 73 307 75 311
rect 99 307 101 311
rect 120 307 122 311
rect 140 307 142 311
rect 145 307 147 311
rect 163 307 165 311
rect 213 307 215 311
rect 218 307 220 311
rect 318 307 320 311
rect 323 307 325 311
rect 213 230 215 234
rect 218 230 220 234
rect 268 234 270 238
rect 294 230 296 234
rect 299 230 301 234
rect 358 234 360 238
rect 384 230 386 234
rect 389 230 391 234
rect 241 226 243 230
rect 13 221 15 225
rect 29 221 31 225
rect 45 221 47 225
rect 68 221 70 225
rect 73 221 75 225
rect 99 221 101 225
rect 120 221 122 225
rect 140 221 142 225
rect 145 221 147 225
rect 163 221 165 225
rect 322 226 324 230
rect 412 226 414 230
rect 13 175 15 179
rect 29 175 31 179
rect 45 175 47 179
rect 68 175 70 179
rect 73 175 75 179
rect 99 175 101 179
rect 120 175 122 179
rect 140 175 142 179
rect 145 175 147 179
rect 163 175 165 179
rect 213 172 215 176
rect 218 172 220 176
rect 294 172 296 176
rect 299 172 301 176
rect 384 172 386 176
rect 389 172 391 176
rect 213 98 215 102
rect 218 98 220 102
rect 241 94 243 98
rect 13 89 15 93
rect 29 89 31 93
rect 45 89 47 93
rect 68 89 70 93
rect 73 89 75 93
rect 99 89 101 93
rect 120 89 122 93
rect 140 89 142 93
rect 145 89 147 93
rect 163 89 165 93
rect 13 43 15 47
rect 29 43 31 47
rect 45 43 47 47
rect 68 43 70 47
rect 73 43 75 47
rect 99 43 101 47
rect 120 43 122 47
rect 140 43 142 47
rect 145 43 147 47
rect 163 43 165 47
rect 247 43 249 47
rect 265 43 267 47
rect 290 43 292 47
rect 306 43 308 47
rect 329 43 331 47
rect 334 43 336 47
rect 360 43 362 47
rect 381 43 383 47
rect 401 43 403 47
rect 406 43 408 47
rect 424 43 426 47
rect 213 36 215 40
rect 218 36 220 40
<< ptransistor >>
rect 8 587 10 595
rect 13 587 15 595
rect 29 587 31 595
rect 45 587 47 595
rect 50 587 52 595
rect 71 587 73 595
rect 87 587 89 595
rect 103 587 105 595
rect 108 587 110 595
rect 124 587 126 595
rect 140 587 142 595
rect 145 587 147 595
rect 161 587 163 595
rect 177 587 179 595
rect 182 587 184 595
rect 203 587 205 595
rect 219 587 221 595
rect 235 587 237 595
rect 240 587 242 595
rect 256 587 258 595
rect 272 587 274 595
rect 277 587 279 595
rect 293 587 295 595
rect 309 587 311 595
rect 314 587 316 595
rect 335 587 337 595
rect 351 587 353 595
rect 367 587 369 595
rect 372 587 374 595
rect 388 587 390 595
rect 404 587 406 595
rect 409 587 411 595
rect 425 587 427 595
rect 441 587 443 595
rect 446 587 448 595
rect 467 587 469 595
rect 483 587 485 595
rect 499 587 501 595
rect 504 587 506 595
rect 520 587 522 595
rect 187 516 189 524
rect 13 503 15 511
rect 29 503 31 511
rect 45 503 47 511
rect 68 503 70 511
rect 73 503 75 511
rect 99 503 101 511
rect 120 503 122 511
rect 140 503 142 511
rect 145 503 147 511
rect 163 503 165 511
rect 213 510 215 518
rect 218 510 220 518
rect 241 516 243 524
rect 268 516 270 524
rect 294 510 296 518
rect 299 510 301 518
rect 322 516 324 524
rect 13 417 15 425
rect 29 417 31 425
rect 45 417 47 425
rect 68 417 70 425
rect 73 417 75 425
rect 99 417 101 425
rect 120 417 122 425
rect 140 417 142 425
rect 145 417 147 425
rect 163 417 165 425
rect 213 418 215 426
rect 218 418 220 426
rect 294 418 296 426
rect 299 418 301 426
rect 13 371 15 379
rect 29 371 31 379
rect 45 371 47 379
rect 68 371 70 379
rect 73 371 75 379
rect 99 371 101 379
rect 120 371 122 379
rect 140 371 142 379
rect 145 371 147 379
rect 163 371 165 379
rect 213 378 215 386
rect 218 378 220 386
rect 241 384 243 392
rect 292 384 294 392
rect 318 378 320 386
rect 323 378 325 386
rect 346 384 348 392
rect 13 285 15 293
rect 29 285 31 293
rect 45 285 47 293
rect 68 285 70 293
rect 73 285 75 293
rect 99 285 101 293
rect 120 285 122 293
rect 140 285 142 293
rect 145 285 147 293
rect 163 285 165 293
rect 213 287 215 295
rect 218 287 220 295
rect 318 287 320 295
rect 323 287 325 295
rect 13 239 15 247
rect 29 239 31 247
rect 45 239 47 247
rect 68 239 70 247
rect 73 239 75 247
rect 99 239 101 247
rect 120 239 122 247
rect 140 239 142 247
rect 145 239 147 247
rect 163 239 165 247
rect 213 246 215 254
rect 218 246 220 254
rect 241 252 243 260
rect 268 252 270 260
rect 294 246 296 254
rect 299 246 301 254
rect 322 252 324 260
rect 358 252 360 260
rect 384 246 386 254
rect 389 246 391 254
rect 412 252 414 260
rect 13 153 15 161
rect 29 153 31 161
rect 45 153 47 161
rect 68 153 70 161
rect 73 153 75 161
rect 99 153 101 161
rect 120 153 122 161
rect 140 153 142 161
rect 145 153 147 161
rect 163 153 165 161
rect 213 152 215 160
rect 218 152 220 160
rect 294 152 296 160
rect 299 152 301 160
rect 384 152 386 160
rect 389 152 391 160
rect 13 107 15 115
rect 29 107 31 115
rect 45 107 47 115
rect 68 107 70 115
rect 73 107 75 115
rect 99 107 101 115
rect 120 107 122 115
rect 140 107 142 115
rect 145 107 147 115
rect 163 107 165 115
rect 213 114 215 122
rect 218 114 220 122
rect 241 120 243 128
rect 13 21 15 29
rect 29 21 31 29
rect 45 21 47 29
rect 68 21 70 29
rect 73 21 75 29
rect 99 21 101 29
rect 120 21 122 29
rect 140 21 142 29
rect 145 21 147 29
rect 163 21 165 29
rect 213 16 215 24
rect 218 16 220 24
rect 247 21 249 29
rect 265 21 267 29
rect 290 21 292 29
rect 306 21 308 29
rect 329 21 331 29
rect 334 21 336 29
rect 360 21 362 29
rect 381 21 383 29
rect 401 21 403 29
rect 406 21 408 29
rect 424 21 426 29
<< ndiffusion >>
rect 7 564 8 568
rect 10 564 13 568
rect 15 564 16 568
rect 28 564 29 568
rect 31 564 32 568
rect 44 564 45 568
rect 47 564 50 568
rect 52 564 53 568
rect 70 564 71 568
rect 73 564 74 568
rect 86 564 87 568
rect 89 564 90 568
rect 102 564 103 568
rect 105 564 108 568
rect 110 564 111 568
rect 123 564 124 568
rect 126 564 127 568
rect 139 564 140 568
rect 142 564 145 568
rect 147 564 148 568
rect 160 564 161 568
rect 163 564 164 568
rect 176 564 177 568
rect 179 564 182 568
rect 184 564 185 568
rect 202 564 203 568
rect 205 564 206 568
rect 218 564 219 568
rect 221 564 222 568
rect 234 564 235 568
rect 237 564 240 568
rect 242 564 243 568
rect 255 564 256 568
rect 258 564 259 568
rect 271 564 272 568
rect 274 564 277 568
rect 279 564 280 568
rect 292 564 293 568
rect 295 564 296 568
rect 308 564 309 568
rect 311 564 314 568
rect 316 564 317 568
rect 334 564 335 568
rect 337 564 338 568
rect 350 564 351 568
rect 353 564 354 568
rect 366 564 367 568
rect 369 564 372 568
rect 374 564 375 568
rect 387 564 388 568
rect 390 564 391 568
rect 403 564 404 568
rect 406 564 409 568
rect 411 564 412 568
rect 424 564 425 568
rect 427 564 428 568
rect 440 564 441 568
rect 443 564 446 568
rect 448 564 449 568
rect 466 564 467 568
rect 469 564 470 568
rect 482 564 483 568
rect 485 564 486 568
rect 498 564 499 568
rect 501 564 504 568
rect 506 564 507 568
rect 519 564 520 568
rect 522 564 523 568
rect 186 498 187 502
rect 189 498 190 502
rect 210 494 213 498
rect 215 494 218 498
rect 220 494 221 498
rect 267 498 268 502
rect 270 498 271 502
rect 291 494 294 498
rect 296 494 299 498
rect 301 494 302 498
rect 240 490 241 494
rect 243 490 244 494
rect 12 485 13 489
rect 15 485 16 489
rect 28 485 29 489
rect 31 485 32 489
rect 44 485 45 489
rect 47 485 48 489
rect 63 485 68 489
rect 70 485 73 489
rect 75 485 76 489
rect 97 485 99 489
rect 101 485 102 489
rect 119 485 120 489
rect 122 485 123 489
rect 135 485 140 489
rect 142 485 145 489
rect 147 485 148 489
rect 162 485 163 489
rect 165 485 166 489
rect 321 490 322 494
rect 324 490 325 494
rect 12 439 13 443
rect 15 439 16 443
rect 28 439 29 443
rect 31 439 32 443
rect 44 439 45 443
rect 47 439 48 443
rect 63 439 68 443
rect 70 439 73 443
rect 75 439 76 443
rect 97 439 99 443
rect 101 439 102 443
rect 119 439 120 443
rect 122 439 123 443
rect 135 439 140 443
rect 142 439 145 443
rect 147 439 148 443
rect 162 439 163 443
rect 165 439 166 443
rect 210 438 213 442
rect 215 438 218 442
rect 220 438 221 442
rect 291 438 294 442
rect 296 438 299 442
rect 301 438 302 442
rect 210 362 213 366
rect 215 362 218 366
rect 220 362 221 366
rect 291 366 292 370
rect 294 366 295 370
rect 315 362 318 366
rect 320 362 323 366
rect 325 362 326 366
rect 240 358 241 362
rect 243 358 244 362
rect 12 353 13 357
rect 15 353 16 357
rect 28 353 29 357
rect 31 353 32 357
rect 44 353 45 357
rect 47 353 48 357
rect 63 353 68 357
rect 70 353 73 357
rect 75 353 76 357
rect 97 353 99 357
rect 101 353 102 357
rect 119 353 120 357
rect 122 353 123 357
rect 135 353 140 357
rect 142 353 145 357
rect 147 353 148 357
rect 162 353 163 357
rect 165 353 166 357
rect 345 358 346 362
rect 348 358 349 362
rect 12 307 13 311
rect 15 307 16 311
rect 28 307 29 311
rect 31 307 32 311
rect 44 307 45 311
rect 47 307 48 311
rect 63 307 68 311
rect 70 307 73 311
rect 75 307 76 311
rect 97 307 99 311
rect 101 307 102 311
rect 119 307 120 311
rect 122 307 123 311
rect 135 307 140 311
rect 142 307 145 311
rect 147 307 148 311
rect 162 307 163 311
rect 165 307 166 311
rect 210 307 213 311
rect 215 307 218 311
rect 220 307 221 311
rect 315 307 318 311
rect 320 307 323 311
rect 325 307 326 311
rect 210 230 213 234
rect 215 230 218 234
rect 220 230 221 234
rect 267 234 268 238
rect 270 234 271 238
rect 291 230 294 234
rect 296 230 299 234
rect 301 230 302 234
rect 357 234 358 238
rect 360 234 361 238
rect 381 230 384 234
rect 386 230 389 234
rect 391 230 392 234
rect 240 226 241 230
rect 243 226 244 230
rect 12 221 13 225
rect 15 221 16 225
rect 28 221 29 225
rect 31 221 32 225
rect 44 221 45 225
rect 47 221 48 225
rect 63 221 68 225
rect 70 221 73 225
rect 75 221 76 225
rect 97 221 99 225
rect 101 221 102 225
rect 119 221 120 225
rect 122 221 123 225
rect 135 221 140 225
rect 142 221 145 225
rect 147 221 148 225
rect 162 221 163 225
rect 165 221 166 225
rect 321 226 322 230
rect 324 226 325 230
rect 411 226 412 230
rect 414 226 415 230
rect 12 175 13 179
rect 15 175 16 179
rect 28 175 29 179
rect 31 175 32 179
rect 44 175 45 179
rect 47 175 48 179
rect 63 175 68 179
rect 70 175 73 179
rect 75 175 76 179
rect 97 175 99 179
rect 101 175 102 179
rect 119 175 120 179
rect 122 175 123 179
rect 135 175 140 179
rect 142 175 145 179
rect 147 175 148 179
rect 162 175 163 179
rect 165 175 166 179
rect 210 172 213 176
rect 215 172 218 176
rect 220 172 221 176
rect 291 172 294 176
rect 296 172 299 176
rect 301 172 302 176
rect 381 172 384 176
rect 386 172 389 176
rect 391 172 392 176
rect 210 98 213 102
rect 215 98 218 102
rect 220 98 221 102
rect 240 94 241 98
rect 243 94 244 98
rect 12 89 13 93
rect 15 89 16 93
rect 28 89 29 93
rect 31 89 32 93
rect 44 89 45 93
rect 47 89 48 93
rect 63 89 68 93
rect 70 89 73 93
rect 75 89 76 93
rect 97 89 99 93
rect 101 89 102 93
rect 119 89 120 93
rect 122 89 123 93
rect 135 89 140 93
rect 142 89 145 93
rect 147 89 148 93
rect 162 89 163 93
rect 165 89 166 93
rect 12 43 13 47
rect 15 43 16 47
rect 28 43 29 47
rect 31 43 32 47
rect 44 43 45 47
rect 47 43 48 47
rect 63 43 68 47
rect 70 43 73 47
rect 75 43 76 47
rect 97 43 99 47
rect 101 43 102 47
rect 119 43 120 47
rect 122 43 123 47
rect 135 43 140 47
rect 142 43 145 47
rect 147 43 148 47
rect 162 43 163 47
rect 165 43 166 47
rect 246 43 247 47
rect 249 43 250 47
rect 254 43 260 47
rect 264 43 265 47
rect 267 43 268 47
rect 289 43 290 47
rect 292 43 293 47
rect 305 43 306 47
rect 308 43 309 47
rect 324 43 329 47
rect 331 43 334 47
rect 336 43 337 47
rect 358 43 360 47
rect 362 43 363 47
rect 380 43 381 47
rect 383 43 384 47
rect 396 43 401 47
rect 403 43 406 47
rect 408 43 409 47
rect 423 43 424 47
rect 426 43 427 47
rect 210 36 213 40
rect 215 36 218 40
rect 220 36 221 40
<< pdiffusion >>
rect 7 587 8 595
rect 10 587 13 595
rect 15 587 16 595
rect 28 587 29 595
rect 31 591 32 595
rect 31 587 36 591
rect 44 587 45 595
rect 47 587 50 595
rect 52 587 53 595
rect 70 587 71 595
rect 73 587 74 595
rect 86 587 87 595
rect 89 591 90 595
rect 89 587 94 591
rect 102 587 103 595
rect 105 587 108 595
rect 110 587 111 595
rect 123 587 124 595
rect 126 587 127 595
rect 139 587 140 595
rect 142 587 145 595
rect 147 587 148 595
rect 160 587 161 595
rect 163 591 164 595
rect 163 587 168 591
rect 176 587 177 595
rect 179 587 182 595
rect 184 587 185 595
rect 202 587 203 595
rect 205 587 206 595
rect 218 587 219 595
rect 221 591 222 595
rect 221 587 226 591
rect 234 587 235 595
rect 237 587 240 595
rect 242 587 243 595
rect 255 587 256 595
rect 258 587 259 595
rect 271 587 272 595
rect 274 587 277 595
rect 279 587 280 595
rect 292 587 293 595
rect 295 591 296 595
rect 295 587 300 591
rect 308 587 309 595
rect 311 587 314 595
rect 316 587 317 595
rect 334 587 335 595
rect 337 587 338 595
rect 350 587 351 595
rect 353 591 354 595
rect 353 587 358 591
rect 366 587 367 595
rect 369 587 372 595
rect 374 587 375 595
rect 387 587 388 595
rect 390 587 391 595
rect 403 587 404 595
rect 406 587 409 595
rect 411 587 412 595
rect 424 587 425 595
rect 427 591 428 595
rect 427 587 432 591
rect 440 587 441 595
rect 443 587 446 595
rect 448 587 449 595
rect 466 587 467 595
rect 469 587 470 595
rect 482 587 483 595
rect 485 591 486 595
rect 485 587 490 591
rect 498 587 499 595
rect 501 587 504 595
rect 506 587 507 595
rect 519 587 520 595
rect 522 587 523 595
rect 186 516 187 524
rect 189 516 190 524
rect 12 503 13 511
rect 15 503 16 511
rect 28 503 29 511
rect 31 503 32 511
rect 44 503 45 511
rect 47 503 48 511
rect 63 503 68 511
rect 70 503 73 511
rect 75 503 76 511
rect 97 503 99 511
rect 101 503 102 511
rect 119 503 120 511
rect 122 503 123 511
rect 135 503 140 511
rect 142 503 145 511
rect 147 503 148 511
rect 162 503 163 511
rect 165 503 166 511
rect 210 510 213 518
rect 215 510 218 518
rect 220 510 221 518
rect 240 516 241 524
rect 243 516 244 524
rect 267 516 268 524
rect 270 516 271 524
rect 291 510 294 518
rect 296 510 299 518
rect 301 510 302 518
rect 321 516 322 524
rect 324 516 325 524
rect 12 417 13 425
rect 15 417 16 425
rect 28 417 29 425
rect 31 417 32 425
rect 44 417 45 425
rect 47 417 48 425
rect 63 417 68 425
rect 70 417 73 425
rect 75 417 76 425
rect 97 417 99 425
rect 101 417 102 425
rect 119 417 120 425
rect 122 417 123 425
rect 135 417 140 425
rect 142 417 145 425
rect 147 417 148 425
rect 162 417 163 425
rect 165 417 166 425
rect 210 418 213 426
rect 215 418 218 426
rect 220 418 221 426
rect 291 418 294 426
rect 296 418 299 426
rect 301 418 302 426
rect 12 371 13 379
rect 15 371 16 379
rect 28 371 29 379
rect 31 371 32 379
rect 44 371 45 379
rect 47 371 48 379
rect 63 371 68 379
rect 70 371 73 379
rect 75 371 76 379
rect 97 371 99 379
rect 101 371 102 379
rect 119 371 120 379
rect 122 371 123 379
rect 135 371 140 379
rect 142 371 145 379
rect 147 371 148 379
rect 162 371 163 379
rect 165 371 166 379
rect 210 378 213 386
rect 215 378 218 386
rect 220 378 221 386
rect 240 384 241 392
rect 243 384 244 392
rect 291 384 292 392
rect 294 384 295 392
rect 315 378 318 386
rect 320 378 323 386
rect 325 378 326 386
rect 345 384 346 392
rect 348 384 349 392
rect 12 285 13 293
rect 15 285 16 293
rect 28 285 29 293
rect 31 285 32 293
rect 44 285 45 293
rect 47 285 48 293
rect 63 285 68 293
rect 70 285 73 293
rect 75 285 76 293
rect 97 285 99 293
rect 101 285 102 293
rect 119 285 120 293
rect 122 285 123 293
rect 135 285 140 293
rect 142 285 145 293
rect 147 285 148 293
rect 162 285 163 293
rect 165 285 166 293
rect 210 287 213 295
rect 215 287 218 295
rect 220 287 221 295
rect 315 287 318 295
rect 320 287 323 295
rect 325 287 326 295
rect 12 239 13 247
rect 15 239 16 247
rect 28 239 29 247
rect 31 239 32 247
rect 44 239 45 247
rect 47 239 48 247
rect 63 239 68 247
rect 70 239 73 247
rect 75 239 76 247
rect 97 239 99 247
rect 101 239 102 247
rect 119 239 120 247
rect 122 239 123 247
rect 135 239 140 247
rect 142 239 145 247
rect 147 239 148 247
rect 162 239 163 247
rect 165 239 166 247
rect 210 246 213 254
rect 215 246 218 254
rect 220 246 221 254
rect 240 252 241 260
rect 243 252 244 260
rect 267 252 268 260
rect 270 252 271 260
rect 291 246 294 254
rect 296 246 299 254
rect 301 246 302 254
rect 321 252 322 260
rect 324 252 325 260
rect 357 252 358 260
rect 360 252 361 260
rect 381 246 384 254
rect 386 246 389 254
rect 391 246 392 254
rect 411 252 412 260
rect 414 252 415 260
rect 12 153 13 161
rect 15 153 16 161
rect 28 153 29 161
rect 31 153 32 161
rect 44 153 45 161
rect 47 153 48 161
rect 63 153 68 161
rect 70 153 73 161
rect 75 153 76 161
rect 97 153 99 161
rect 101 153 102 161
rect 119 153 120 161
rect 122 153 123 161
rect 135 153 140 161
rect 142 153 145 161
rect 147 153 148 161
rect 162 153 163 161
rect 165 153 166 161
rect 210 152 213 160
rect 215 152 218 160
rect 220 152 221 160
rect 291 152 294 160
rect 296 152 299 160
rect 301 152 302 160
rect 381 152 384 160
rect 386 152 389 160
rect 391 152 392 160
rect 12 107 13 115
rect 15 107 16 115
rect 28 107 29 115
rect 31 107 32 115
rect 44 107 45 115
rect 47 107 48 115
rect 63 107 68 115
rect 70 107 73 115
rect 75 107 76 115
rect 97 107 99 115
rect 101 107 102 115
rect 119 107 120 115
rect 122 107 123 115
rect 135 107 140 115
rect 142 107 145 115
rect 147 107 148 115
rect 162 107 163 115
rect 165 107 166 115
rect 210 114 213 122
rect 215 114 218 122
rect 220 114 221 122
rect 240 120 241 128
rect 243 120 244 128
rect 12 21 13 29
rect 15 21 16 29
rect 28 21 29 29
rect 31 21 32 29
rect 44 21 45 29
rect 47 21 48 29
rect 63 21 68 29
rect 70 21 73 29
rect 75 21 76 29
rect 97 21 99 29
rect 101 21 102 29
rect 119 21 120 29
rect 122 21 123 29
rect 135 21 140 29
rect 142 21 145 29
rect 147 21 148 29
rect 162 21 163 29
rect 165 21 166 29
rect 210 16 213 24
rect 215 16 218 24
rect 220 16 221 24
rect 246 21 247 29
rect 249 21 250 29
rect 254 21 260 29
rect 264 21 265 29
rect 267 21 268 29
rect 289 21 290 29
rect 292 21 293 29
rect 305 21 306 29
rect 308 21 309 29
rect 324 21 329 29
rect 331 21 334 29
rect 336 21 337 29
rect 358 21 360 29
rect 362 21 363 29
rect 380 21 381 29
rect 383 21 384 29
rect 396 21 401 29
rect 403 21 406 29
rect 408 21 409 29
rect 423 21 424 29
rect 426 21 427 29
<< ndcontact >>
rect 3 564 7 568
rect 16 564 20 568
rect 24 564 28 568
rect 32 564 36 568
rect 40 564 44 568
rect 53 564 57 568
rect 66 564 70 568
rect 74 564 78 568
rect 82 564 86 568
rect 90 564 94 568
rect 98 564 102 568
rect 111 564 115 568
rect 119 564 123 568
rect 127 564 131 568
rect 135 564 139 568
rect 148 564 152 568
rect 156 564 160 568
rect 164 564 168 568
rect 172 564 176 568
rect 185 564 189 568
rect 198 564 202 568
rect 206 564 210 568
rect 214 564 218 568
rect 222 564 226 568
rect 230 564 234 568
rect 243 564 247 568
rect 251 564 255 568
rect 259 564 263 568
rect 267 564 271 568
rect 280 564 284 568
rect 288 564 292 568
rect 296 564 300 568
rect 304 564 308 568
rect 317 564 321 568
rect 330 564 334 568
rect 338 564 342 568
rect 346 564 350 568
rect 354 564 358 568
rect 362 564 366 568
rect 375 564 379 568
rect 383 564 387 568
rect 391 564 395 568
rect 399 564 403 568
rect 412 564 416 568
rect 420 564 424 568
rect 428 564 432 568
rect 436 564 440 568
rect 449 564 453 568
rect 462 564 466 568
rect 470 564 474 568
rect 478 564 482 568
rect 486 564 490 568
rect 494 564 498 568
rect 507 564 511 568
rect 515 564 519 568
rect 523 564 527 568
rect 182 498 186 502
rect 190 498 194 502
rect 206 494 210 498
rect 221 494 225 498
rect 263 498 267 502
rect 271 498 275 502
rect 287 494 291 498
rect 302 494 306 498
rect 236 490 240 494
rect 244 490 248 494
rect 8 485 12 489
rect 16 485 20 489
rect 24 485 28 489
rect 32 485 36 489
rect 40 485 44 489
rect 48 485 52 489
rect 59 485 63 489
rect 76 485 80 489
rect 93 485 97 489
rect 102 485 106 489
rect 115 485 119 489
rect 123 485 127 489
rect 131 485 135 489
rect 148 485 152 489
rect 158 485 162 489
rect 166 485 170 489
rect 317 490 321 494
rect 325 490 329 494
rect 8 439 12 443
rect 16 439 20 443
rect 24 439 28 443
rect 32 439 36 443
rect 40 439 44 443
rect 48 439 52 443
rect 59 439 63 443
rect 76 439 80 443
rect 93 439 97 443
rect 102 439 106 443
rect 115 439 119 443
rect 123 439 127 443
rect 131 439 135 443
rect 148 439 152 443
rect 158 439 162 443
rect 166 439 170 443
rect 206 438 210 442
rect 221 438 225 442
rect 287 438 291 442
rect 302 438 306 442
rect 206 362 210 366
rect 221 362 225 366
rect 287 366 291 370
rect 295 366 299 370
rect 311 362 315 366
rect 326 362 330 366
rect 236 358 240 362
rect 244 358 248 362
rect 8 353 12 357
rect 16 353 20 357
rect 24 353 28 357
rect 32 353 36 357
rect 40 353 44 357
rect 48 353 52 357
rect 59 353 63 357
rect 76 353 80 357
rect 93 353 97 357
rect 102 353 106 357
rect 115 353 119 357
rect 123 353 127 357
rect 131 353 135 357
rect 148 353 152 357
rect 158 353 162 357
rect 166 353 170 357
rect 341 358 345 362
rect 349 358 353 362
rect 8 307 12 311
rect 16 307 20 311
rect 24 307 28 311
rect 32 307 36 311
rect 40 307 44 311
rect 48 307 52 311
rect 59 307 63 311
rect 76 307 80 311
rect 93 307 97 311
rect 102 307 106 311
rect 115 307 119 311
rect 123 307 127 311
rect 131 307 135 311
rect 148 307 152 311
rect 158 307 162 311
rect 166 307 170 311
rect 206 307 210 311
rect 221 307 225 311
rect 311 307 315 311
rect 326 307 330 311
rect 206 230 210 234
rect 221 230 225 234
rect 263 234 267 238
rect 271 234 275 238
rect 287 230 291 234
rect 302 230 306 234
rect 353 234 357 238
rect 361 234 365 238
rect 377 230 381 234
rect 392 230 396 234
rect 236 226 240 230
rect 244 226 248 230
rect 8 221 12 225
rect 16 221 20 225
rect 24 221 28 225
rect 32 221 36 225
rect 40 221 44 225
rect 48 221 52 225
rect 59 221 63 225
rect 76 221 80 225
rect 93 221 97 225
rect 102 221 106 225
rect 115 221 119 225
rect 123 221 127 225
rect 131 221 135 225
rect 148 221 152 225
rect 158 221 162 225
rect 166 221 170 225
rect 317 226 321 230
rect 325 226 329 230
rect 407 226 411 230
rect 415 226 419 230
rect 8 175 12 179
rect 16 175 20 179
rect 24 175 28 179
rect 32 175 36 179
rect 40 175 44 179
rect 48 175 52 179
rect 59 175 63 179
rect 76 175 80 179
rect 93 175 97 179
rect 102 175 106 179
rect 115 175 119 179
rect 123 175 127 179
rect 131 175 135 179
rect 148 175 152 179
rect 158 175 162 179
rect 166 175 170 179
rect 206 172 210 176
rect 221 172 225 176
rect 287 172 291 176
rect 302 172 306 176
rect 377 172 381 176
rect 392 172 396 176
rect 206 98 210 102
rect 221 98 225 102
rect 236 94 240 98
rect 244 94 248 98
rect 8 89 12 93
rect 16 89 20 93
rect 24 89 28 93
rect 32 89 36 93
rect 40 89 44 93
rect 48 89 52 93
rect 59 89 63 93
rect 76 89 80 93
rect 93 89 97 93
rect 102 89 106 93
rect 115 89 119 93
rect 123 89 127 93
rect 131 89 135 93
rect 148 89 152 93
rect 158 89 162 93
rect 166 89 170 93
rect 8 43 12 47
rect 16 43 20 47
rect 24 43 28 47
rect 32 43 36 47
rect 40 43 44 47
rect 48 43 52 47
rect 59 43 63 47
rect 76 43 80 47
rect 93 43 97 47
rect 102 43 106 47
rect 115 43 119 47
rect 123 43 127 47
rect 131 43 135 47
rect 148 43 152 47
rect 158 43 162 47
rect 166 43 170 47
rect 242 43 246 47
rect 250 43 254 47
rect 260 43 264 47
rect 268 43 272 47
rect 277 43 281 47
rect 285 43 289 47
rect 293 43 297 47
rect 301 43 305 47
rect 309 43 313 47
rect 320 43 324 47
rect 337 43 341 47
rect 354 43 358 47
rect 363 43 367 47
rect 376 43 380 47
rect 384 43 388 47
rect 392 43 396 47
rect 409 43 413 47
rect 419 43 423 47
rect 427 43 431 47
rect 206 36 210 40
rect 221 36 225 40
<< pdcontact >>
rect 3 587 7 595
rect 16 587 20 595
rect 24 587 28 595
rect 32 591 36 595
rect 40 587 44 595
rect 53 587 57 595
rect 66 587 70 595
rect 74 587 78 595
rect 82 587 86 595
rect 90 591 94 595
rect 98 587 102 595
rect 111 587 115 595
rect 119 587 123 595
rect 127 587 131 595
rect 135 587 139 595
rect 148 587 152 595
rect 156 587 160 595
rect 164 591 168 595
rect 172 587 176 595
rect 185 587 189 595
rect 198 587 202 595
rect 206 587 210 595
rect 214 587 218 595
rect 222 591 226 595
rect 230 587 234 595
rect 243 587 247 595
rect 251 587 255 595
rect 259 587 263 595
rect 267 587 271 595
rect 280 587 284 595
rect 288 587 292 595
rect 296 591 300 595
rect 304 587 308 595
rect 317 587 321 595
rect 330 587 334 595
rect 338 587 342 595
rect 346 587 350 595
rect 354 591 358 595
rect 362 587 366 595
rect 375 587 379 595
rect 383 587 387 595
rect 391 587 395 595
rect 399 587 403 595
rect 412 587 416 595
rect 420 587 424 595
rect 428 591 432 595
rect 436 587 440 595
rect 449 587 453 595
rect 462 587 466 595
rect 470 587 474 595
rect 478 587 482 595
rect 486 591 490 595
rect 494 587 498 595
rect 507 587 511 595
rect 515 587 519 595
rect 523 587 527 595
rect 182 516 186 524
rect 190 516 194 524
rect 8 503 12 511
rect 16 503 20 511
rect 24 503 28 511
rect 32 503 36 511
rect 40 503 44 511
rect 48 503 52 511
rect 59 503 63 511
rect 76 503 80 511
rect 93 503 97 511
rect 102 503 106 511
rect 115 503 119 511
rect 123 503 127 511
rect 131 503 135 511
rect 148 503 152 511
rect 158 503 162 511
rect 166 503 170 511
rect 206 510 210 518
rect 221 510 225 518
rect 236 516 240 524
rect 244 516 248 524
rect 263 516 267 524
rect 271 516 275 524
rect 287 510 291 518
rect 302 510 306 518
rect 317 516 321 524
rect 325 516 329 524
rect 8 417 12 425
rect 16 417 20 425
rect 24 417 28 425
rect 32 417 36 425
rect 40 417 44 425
rect 48 417 52 425
rect 59 417 63 425
rect 76 417 80 425
rect 93 417 97 425
rect 102 417 106 425
rect 115 417 119 425
rect 123 417 127 425
rect 131 417 135 425
rect 148 417 152 425
rect 158 417 162 425
rect 166 417 170 425
rect 206 418 210 426
rect 221 418 225 426
rect 287 418 291 426
rect 302 418 306 426
rect 8 371 12 379
rect 16 371 20 379
rect 24 371 28 379
rect 32 371 36 379
rect 40 371 44 379
rect 48 371 52 379
rect 59 371 63 379
rect 76 371 80 379
rect 93 371 97 379
rect 102 371 106 379
rect 115 371 119 379
rect 123 371 127 379
rect 131 371 135 379
rect 148 371 152 379
rect 158 371 162 379
rect 166 371 170 379
rect 206 378 210 386
rect 221 378 225 386
rect 236 384 240 392
rect 244 384 248 392
rect 287 384 291 392
rect 295 384 299 392
rect 311 378 315 386
rect 326 378 330 386
rect 341 384 345 392
rect 349 384 353 392
rect 8 285 12 293
rect 16 285 20 293
rect 24 285 28 293
rect 32 285 36 293
rect 40 285 44 293
rect 48 285 52 293
rect 59 285 63 293
rect 76 285 80 293
rect 93 285 97 293
rect 102 285 106 293
rect 115 285 119 293
rect 123 285 127 293
rect 131 285 135 293
rect 148 285 152 293
rect 158 285 162 293
rect 166 285 170 293
rect 206 287 210 295
rect 221 287 225 295
rect 311 287 315 295
rect 326 287 330 295
rect 8 239 12 247
rect 16 239 20 247
rect 24 239 28 247
rect 32 239 36 247
rect 40 239 44 247
rect 48 239 52 247
rect 59 239 63 247
rect 76 239 80 247
rect 93 239 97 247
rect 102 239 106 247
rect 115 239 119 247
rect 123 239 127 247
rect 131 239 135 247
rect 148 239 152 247
rect 158 239 162 247
rect 166 239 170 247
rect 206 246 210 254
rect 221 246 225 254
rect 236 252 240 260
rect 244 252 248 260
rect 263 252 267 260
rect 271 252 275 260
rect 287 246 291 254
rect 302 246 306 254
rect 317 252 321 260
rect 325 252 329 260
rect 353 252 357 260
rect 361 252 365 260
rect 377 246 381 254
rect 392 246 396 254
rect 407 252 411 260
rect 415 252 419 260
rect 8 153 12 161
rect 16 153 20 161
rect 24 153 28 161
rect 32 153 36 161
rect 40 153 44 161
rect 48 153 52 161
rect 59 153 63 161
rect 76 153 80 161
rect 93 153 97 161
rect 102 153 106 161
rect 115 153 119 161
rect 123 153 127 161
rect 131 153 135 161
rect 148 153 152 161
rect 158 153 162 161
rect 166 153 170 161
rect 206 152 210 160
rect 221 152 225 160
rect 287 152 291 160
rect 302 152 306 160
rect 377 152 381 160
rect 392 152 396 160
rect 8 107 12 115
rect 16 107 20 115
rect 24 107 28 115
rect 32 107 36 115
rect 40 107 44 115
rect 48 107 52 115
rect 59 107 63 115
rect 76 107 80 115
rect 93 107 97 115
rect 102 107 106 115
rect 115 107 119 115
rect 123 107 127 115
rect 131 107 135 115
rect 148 107 152 115
rect 158 107 162 115
rect 166 107 170 115
rect 206 114 210 122
rect 221 114 225 122
rect 236 120 240 128
rect 244 120 248 128
rect 8 21 12 29
rect 16 21 20 29
rect 24 21 28 29
rect 32 21 36 29
rect 40 21 44 29
rect 48 21 52 29
rect 59 21 63 29
rect 76 21 80 29
rect 93 21 97 29
rect 102 21 106 29
rect 115 21 119 29
rect 123 21 127 29
rect 131 21 135 29
rect 148 21 152 29
rect 158 21 162 29
rect 166 21 170 29
rect 206 16 210 24
rect 221 16 225 24
rect 242 21 246 29
rect 250 21 254 29
rect 260 21 264 29
rect 268 21 272 29
rect 277 21 281 29
rect 285 21 289 29
rect 293 21 297 29
rect 301 21 305 29
rect 309 21 313 29
rect 320 21 324 29
rect 337 21 341 29
rect 354 21 358 29
rect 363 21 367 29
rect 376 21 380 29
rect 384 21 388 29
rect 392 21 396 29
rect 409 21 413 29
rect 419 21 423 29
rect 427 21 431 29
<< psubstratepcontact >>
rect 33 548 37 552
rect 61 548 65 552
rect 91 548 95 552
rect 165 548 169 552
rect 193 548 197 552
rect 223 548 227 552
rect 297 548 301 552
rect 325 548 329 552
rect 355 548 359 552
rect 429 548 433 552
rect 457 548 461 552
rect 487 548 491 552
rect 14 462 18 466
rect 49 462 53 466
rect 175 462 179 466
rect 199 462 203 466
rect 253 462 260 466
rect 280 462 284 466
rect 334 462 338 466
rect 14 330 18 334
rect 49 330 53 334
rect 175 330 179 334
rect 199 330 203 334
rect 253 330 257 334
rect 280 330 284 334
rect 304 330 308 334
rect 14 198 18 202
rect 49 198 53 202
rect 175 198 179 202
rect 199 198 203 202
rect 253 198 260 202
rect 280 198 284 202
rect 334 198 338 202
rect 370 198 374 202
rect 424 198 428 202
rect 14 66 18 70
rect 49 66 53 70
rect 175 66 179 70
rect 199 66 203 70
rect 310 66 314 70
<< nsubstratencontact >>
rect 33 605 37 609
rect 61 605 65 609
rect 91 605 95 609
rect 128 605 132 609
rect 165 605 169 609
rect 193 605 197 609
rect 223 605 227 609
rect 260 605 264 609
rect 297 605 301 609
rect 325 605 329 609
rect 355 605 359 609
rect 392 605 396 609
rect 429 605 433 609
rect 457 605 461 609
rect 487 605 491 609
rect 524 605 528 609
rect 23 528 27 532
rect 52 528 56 532
rect 77 528 81 532
rect 119 528 123 532
rect 175 528 179 532
rect 199 528 203 532
rect 253 528 257 532
rect 280 528 284 532
rect 334 528 338 532
rect 23 396 27 400
rect 52 396 56 400
rect 77 396 81 400
rect 119 396 123 400
rect 175 396 179 400
rect 199 396 203 400
rect 253 396 257 400
rect 280 396 284 400
rect 342 396 346 400
rect 23 264 27 268
rect 52 264 56 268
rect 77 264 81 268
rect 119 264 123 268
rect 175 264 179 268
rect 199 264 203 268
rect 253 264 257 268
rect 280 264 284 268
rect 334 264 338 268
rect 342 264 346 268
rect 370 264 374 268
rect 424 264 428 268
rect 23 132 27 136
rect 52 132 56 136
rect 77 132 81 136
rect 119 132 123 136
rect 175 132 179 136
rect 199 132 203 136
rect 253 132 257 136
rect 280 132 284 136
rect 370 132 374 136
rect 23 0 27 4
rect 52 0 56 4
rect 77 0 81 4
rect 119 0 123 4
rect 199 0 203 4
rect 253 0 257 4
rect 284 0 288 4
rect 313 0 317 4
rect 338 0 342 4
rect 380 0 384 4
<< polysilicon >>
rect 8 595 10 597
rect 13 595 15 598
rect 29 595 31 597
rect 45 595 47 597
rect 50 595 52 598
rect 71 595 73 598
rect 87 595 89 598
rect 103 595 105 597
rect 108 595 110 598
rect 124 595 126 597
rect 140 595 142 597
rect 145 595 147 598
rect 161 595 163 597
rect 177 595 179 597
rect 182 595 184 598
rect 203 595 205 598
rect 219 595 221 598
rect 235 595 237 597
rect 240 595 242 598
rect 256 595 258 597
rect 272 595 274 597
rect 277 595 279 598
rect 293 595 295 597
rect 309 595 311 597
rect 314 595 316 598
rect 335 595 337 598
rect 351 595 353 598
rect 367 595 369 597
rect 372 595 374 598
rect 388 595 390 597
rect 404 595 406 597
rect 409 595 411 598
rect 425 595 427 597
rect 441 595 443 597
rect 446 595 448 598
rect 467 595 469 598
rect 483 595 485 598
rect 499 595 501 597
rect 504 595 506 598
rect 520 595 522 597
rect 8 582 10 587
rect 13 585 15 587
rect 8 568 10 578
rect 13 568 15 575
rect 29 568 31 587
rect 45 578 47 587
rect 50 585 52 587
rect 71 585 73 587
rect 87 584 89 587
rect 45 568 47 571
rect 50 568 52 570
rect 71 568 73 570
rect 87 568 89 580
rect 103 578 105 587
rect 108 585 110 587
rect 124 579 126 587
rect 140 582 142 587
rect 145 585 147 587
rect 103 568 105 571
rect 108 568 110 570
rect 124 568 126 575
rect 140 568 142 578
rect 145 568 147 575
rect 161 568 163 587
rect 177 578 179 587
rect 182 585 184 587
rect 203 585 205 587
rect 219 584 221 587
rect 177 568 179 571
rect 182 568 184 570
rect 203 568 205 570
rect 219 568 221 580
rect 235 578 237 587
rect 240 585 242 587
rect 256 579 258 587
rect 272 582 274 587
rect 277 585 279 587
rect 235 568 237 571
rect 240 568 242 570
rect 256 568 258 575
rect 272 568 274 578
rect 277 568 279 575
rect 293 568 295 587
rect 309 578 311 587
rect 314 585 316 587
rect 335 585 337 587
rect 351 584 353 587
rect 309 568 311 571
rect 314 568 316 570
rect 335 568 337 570
rect 351 568 353 580
rect 367 578 369 587
rect 372 585 374 587
rect 388 579 390 587
rect 404 582 406 587
rect 409 585 411 587
rect 367 568 369 571
rect 372 568 374 570
rect 388 568 390 575
rect 404 568 406 578
rect 409 568 411 575
rect 425 568 427 587
rect 441 578 443 587
rect 446 585 448 587
rect 467 585 469 587
rect 483 584 485 587
rect 441 568 443 571
rect 446 568 448 570
rect 467 568 469 570
rect 483 568 485 580
rect 499 578 501 587
rect 504 585 506 587
rect 520 579 522 587
rect 499 568 501 571
rect 504 568 506 570
rect 520 568 522 575
rect 8 562 10 564
rect 13 561 15 564
rect 29 562 31 564
rect 45 562 47 564
rect 50 559 52 564
rect 71 559 73 564
rect 87 562 89 564
rect 103 562 105 564
rect 108 559 110 564
rect 124 562 126 564
rect 140 562 142 564
rect 145 561 147 564
rect 161 562 163 564
rect 177 562 179 564
rect 182 559 184 564
rect 203 559 205 564
rect 219 562 221 564
rect 235 562 237 564
rect 240 559 242 564
rect 256 562 258 564
rect 272 562 274 564
rect 277 561 279 564
rect 293 562 295 564
rect 309 562 311 564
rect 314 559 316 564
rect 335 559 337 564
rect 351 562 353 564
rect 367 562 369 564
rect 372 559 374 564
rect 388 562 390 564
rect 404 562 406 564
rect 409 561 411 564
rect 425 562 427 564
rect 441 562 443 564
rect 446 559 448 564
rect 467 559 469 564
rect 483 562 485 564
rect 499 562 501 564
rect 504 559 506 564
rect 520 562 522 564
rect 187 524 189 526
rect 29 518 31 521
rect 73 518 75 521
rect 99 518 101 521
rect 145 518 147 521
rect 99 514 100 518
rect 213 518 215 522
rect 241 524 243 526
rect 268 524 270 526
rect 218 518 220 521
rect 13 511 15 513
rect 29 511 31 514
rect 45 511 47 513
rect 68 511 70 513
rect 73 511 75 514
rect 99 511 101 514
rect 120 511 122 514
rect 140 511 142 513
rect 145 511 147 514
rect 163 511 165 513
rect 13 489 15 503
rect 29 501 31 503
rect 29 489 31 491
rect 45 489 47 503
rect 68 498 70 503
rect 73 501 75 503
rect 99 501 101 503
rect 64 494 70 498
rect 68 489 70 494
rect 73 489 75 491
rect 99 489 101 491
rect 120 489 122 503
rect 140 498 142 503
rect 145 501 147 503
rect 136 494 142 498
rect 140 489 142 494
rect 145 489 147 491
rect 163 489 165 503
rect 187 502 189 516
rect 294 518 296 522
rect 322 524 324 526
rect 299 518 301 521
rect 213 507 215 510
rect 218 508 220 510
rect 214 503 215 507
rect 213 498 215 503
rect 218 498 220 500
rect 187 496 189 498
rect 241 494 243 516
rect 268 502 270 516
rect 294 507 296 510
rect 299 508 301 510
rect 295 503 296 507
rect 294 498 296 503
rect 299 498 301 500
rect 268 496 270 498
rect 322 494 324 516
rect 213 492 215 494
rect 218 489 220 494
rect 294 492 296 494
rect 241 488 243 490
rect 299 489 301 494
rect 322 488 324 490
rect 13 483 15 485
rect 29 481 31 485
rect 45 483 47 485
rect 68 483 70 485
rect 30 477 31 481
rect 73 480 75 485
rect 99 481 101 485
rect 120 483 122 485
rect 140 483 142 485
rect 29 474 31 477
rect 74 476 75 480
rect 100 477 101 481
rect 145 480 147 485
rect 163 483 165 485
rect 73 474 75 476
rect 99 473 101 477
rect 146 476 147 480
rect 145 474 147 476
rect 29 451 31 454
rect 73 452 75 454
rect 30 447 31 451
rect 74 448 75 452
rect 99 451 101 455
rect 145 452 147 454
rect 13 443 15 445
rect 29 443 31 447
rect 45 443 47 445
rect 68 443 70 445
rect 73 443 75 448
rect 100 447 101 451
rect 146 448 147 452
rect 99 443 101 447
rect 120 443 122 445
rect 140 443 142 445
rect 145 443 147 448
rect 163 443 165 445
rect 213 442 215 445
rect 218 442 220 445
rect 294 442 296 445
rect 299 442 301 445
rect 13 425 15 439
rect 29 437 31 439
rect 29 425 31 427
rect 45 425 47 439
rect 68 434 70 439
rect 73 437 75 439
rect 99 437 101 439
rect 64 430 70 434
rect 68 425 70 430
rect 73 425 75 427
rect 99 425 101 427
rect 120 425 122 439
rect 140 434 142 439
rect 145 437 147 439
rect 136 430 142 434
rect 140 425 142 430
rect 145 425 147 427
rect 163 425 165 439
rect 213 426 215 438
rect 218 436 220 438
rect 218 426 220 428
rect 294 426 296 438
rect 299 436 301 438
rect 299 426 301 428
rect 13 415 15 417
rect 29 414 31 417
rect 45 415 47 417
rect 68 415 70 417
rect 73 414 75 417
rect 99 414 101 417
rect 120 414 122 417
rect 140 415 142 417
rect 145 414 147 417
rect 163 415 165 417
rect 213 416 215 418
rect 99 410 100 414
rect 218 413 220 418
rect 294 416 296 418
rect 299 413 301 418
rect 29 407 31 410
rect 73 407 75 410
rect 99 407 101 410
rect 145 407 147 410
rect 29 386 31 389
rect 73 386 75 389
rect 99 386 101 389
rect 145 386 147 389
rect 213 386 215 390
rect 241 392 243 394
rect 292 392 294 394
rect 218 386 220 389
rect 99 382 100 386
rect 13 379 15 381
rect 29 379 31 382
rect 45 379 47 381
rect 68 379 70 381
rect 73 379 75 382
rect 99 379 101 382
rect 120 379 122 382
rect 140 379 142 381
rect 145 379 147 382
rect 163 379 165 381
rect 318 386 320 390
rect 346 392 348 394
rect 323 386 325 389
rect 213 375 215 378
rect 218 376 220 378
rect 214 371 215 375
rect 13 357 15 371
rect 29 369 31 371
rect 29 357 31 359
rect 45 357 47 371
rect 68 366 70 371
rect 73 369 75 371
rect 99 369 101 371
rect 64 362 70 366
rect 68 357 70 362
rect 73 357 75 359
rect 99 357 101 359
rect 120 357 122 371
rect 140 366 142 371
rect 145 369 147 371
rect 136 362 142 366
rect 140 357 142 362
rect 145 357 147 359
rect 163 357 165 371
rect 213 366 215 371
rect 218 366 220 368
rect 241 362 243 384
rect 292 370 294 384
rect 318 375 320 378
rect 323 376 325 378
rect 319 371 320 375
rect 318 366 320 371
rect 323 366 325 368
rect 292 364 294 366
rect 346 362 348 384
rect 213 360 215 362
rect 218 357 220 362
rect 318 360 320 362
rect 241 356 243 358
rect 323 357 325 362
rect 346 356 348 358
rect 13 351 15 353
rect 29 349 31 353
rect 45 351 47 353
rect 68 351 70 353
rect 30 345 31 349
rect 73 348 75 353
rect 99 349 101 353
rect 120 351 122 353
rect 140 351 142 353
rect 29 342 31 345
rect 74 344 75 348
rect 100 345 101 349
rect 145 348 147 353
rect 163 351 165 353
rect 73 342 75 344
rect 99 341 101 345
rect 146 344 147 348
rect 145 342 147 344
rect 29 319 31 322
rect 73 320 75 322
rect 30 315 31 319
rect 74 316 75 320
rect 99 319 101 323
rect 145 320 147 322
rect 13 311 15 313
rect 29 311 31 315
rect 45 311 47 313
rect 68 311 70 313
rect 73 311 75 316
rect 100 315 101 319
rect 146 316 147 320
rect 99 311 101 315
rect 120 311 122 313
rect 140 311 142 313
rect 145 311 147 316
rect 163 311 165 313
rect 213 311 215 314
rect 218 311 220 314
rect 318 311 320 314
rect 323 311 325 314
rect 13 293 15 307
rect 29 305 31 307
rect 29 293 31 295
rect 45 293 47 307
rect 68 302 70 307
rect 73 305 75 307
rect 99 305 101 307
rect 64 298 70 302
rect 68 293 70 298
rect 73 293 75 295
rect 99 293 101 295
rect 120 293 122 307
rect 140 302 142 307
rect 145 305 147 307
rect 136 298 142 302
rect 140 293 142 298
rect 145 293 147 295
rect 163 293 165 307
rect 213 295 215 307
rect 218 305 220 307
rect 218 295 220 297
rect 318 295 320 307
rect 323 305 325 307
rect 323 295 325 297
rect 213 285 215 287
rect 13 283 15 285
rect 29 282 31 285
rect 45 283 47 285
rect 68 283 70 285
rect 73 282 75 285
rect 99 282 101 285
rect 120 282 122 285
rect 140 283 142 285
rect 145 282 147 285
rect 163 283 165 285
rect 218 282 220 287
rect 318 285 320 287
rect 323 282 325 287
rect 99 278 100 282
rect 29 275 31 278
rect 73 275 75 278
rect 99 275 101 278
rect 145 275 147 278
rect 29 254 31 257
rect 73 254 75 257
rect 99 254 101 257
rect 145 254 147 257
rect 213 254 215 258
rect 241 260 243 262
rect 268 260 270 262
rect 218 254 220 257
rect 99 250 100 254
rect 13 247 15 249
rect 29 247 31 250
rect 45 247 47 249
rect 68 247 70 249
rect 73 247 75 250
rect 99 247 101 250
rect 120 247 122 250
rect 140 247 142 249
rect 145 247 147 250
rect 163 247 165 249
rect 294 254 296 258
rect 322 260 324 262
rect 358 260 360 262
rect 299 254 301 257
rect 213 243 215 246
rect 218 244 220 246
rect 214 239 215 243
rect 13 225 15 239
rect 29 237 31 239
rect 29 225 31 227
rect 45 225 47 239
rect 68 234 70 239
rect 73 237 75 239
rect 99 237 101 239
rect 64 230 70 234
rect 68 225 70 230
rect 73 225 75 227
rect 99 225 101 227
rect 120 225 122 239
rect 140 234 142 239
rect 145 237 147 239
rect 136 230 142 234
rect 140 225 142 230
rect 145 225 147 227
rect 163 225 165 239
rect 213 234 215 239
rect 218 234 220 236
rect 241 230 243 252
rect 268 238 270 252
rect 384 254 386 258
rect 412 260 414 262
rect 389 254 391 257
rect 294 243 296 246
rect 299 244 301 246
rect 295 239 296 243
rect 294 234 296 239
rect 299 234 301 236
rect 268 232 270 234
rect 322 230 324 252
rect 358 238 360 252
rect 384 243 386 246
rect 389 244 391 246
rect 385 239 386 243
rect 384 234 386 239
rect 389 234 391 236
rect 358 232 360 234
rect 412 230 414 252
rect 213 228 215 230
rect 218 225 220 230
rect 294 228 296 230
rect 241 224 243 226
rect 299 225 301 230
rect 384 228 386 230
rect 322 224 324 226
rect 389 225 391 230
rect 412 224 414 226
rect 13 219 15 221
rect 29 217 31 221
rect 45 219 47 221
rect 68 219 70 221
rect 30 213 31 217
rect 73 216 75 221
rect 99 217 101 221
rect 120 219 122 221
rect 140 219 142 221
rect 29 210 31 213
rect 74 212 75 216
rect 100 213 101 217
rect 145 216 147 221
rect 163 219 165 221
rect 73 210 75 212
rect 99 209 101 213
rect 146 212 147 216
rect 145 210 147 212
rect 29 187 31 190
rect 73 188 75 190
rect 30 183 31 187
rect 74 184 75 188
rect 99 187 101 191
rect 145 188 147 190
rect 13 179 15 181
rect 29 179 31 183
rect 45 179 47 181
rect 68 179 70 181
rect 73 179 75 184
rect 100 183 101 187
rect 146 184 147 188
rect 99 179 101 183
rect 120 179 122 181
rect 140 179 142 181
rect 145 179 147 184
rect 163 179 165 181
rect 213 176 215 179
rect 218 176 220 179
rect 294 176 296 179
rect 299 176 301 179
rect 384 176 386 179
rect 389 176 391 179
rect 13 161 15 175
rect 29 173 31 175
rect 29 161 31 163
rect 45 161 47 175
rect 68 170 70 175
rect 73 173 75 175
rect 99 173 101 175
rect 64 166 70 170
rect 68 161 70 166
rect 73 161 75 163
rect 99 161 101 163
rect 120 161 122 175
rect 140 170 142 175
rect 145 173 147 175
rect 136 166 142 170
rect 140 161 142 166
rect 145 161 147 163
rect 163 161 165 175
rect 213 160 215 172
rect 218 170 220 172
rect 218 160 220 162
rect 294 160 296 172
rect 299 170 301 172
rect 299 160 301 162
rect 384 160 386 172
rect 389 170 391 172
rect 389 160 391 162
rect 13 151 15 153
rect 29 150 31 153
rect 45 151 47 153
rect 68 151 70 153
rect 73 150 75 153
rect 99 150 101 153
rect 120 150 122 153
rect 140 151 142 153
rect 145 150 147 153
rect 163 151 165 153
rect 213 150 215 152
rect 99 146 100 150
rect 218 147 220 152
rect 294 150 296 152
rect 299 147 301 152
rect 384 150 386 152
rect 389 147 391 152
rect 29 143 31 146
rect 73 143 75 146
rect 99 143 101 146
rect 145 143 147 146
rect 29 122 31 125
rect 73 122 75 125
rect 99 122 101 125
rect 145 122 147 125
rect 213 122 215 126
rect 241 128 243 130
rect 218 122 220 125
rect 99 118 100 122
rect 13 115 15 117
rect 29 115 31 118
rect 45 115 47 117
rect 68 115 70 117
rect 73 115 75 118
rect 99 115 101 118
rect 120 115 122 118
rect 140 115 142 117
rect 145 115 147 118
rect 163 115 165 117
rect 213 111 215 114
rect 218 112 220 114
rect 214 107 215 111
rect 13 93 15 107
rect 29 105 31 107
rect 29 93 31 95
rect 45 93 47 107
rect 68 102 70 107
rect 73 105 75 107
rect 99 105 101 107
rect 64 98 70 102
rect 68 93 70 98
rect 73 93 75 95
rect 99 93 101 95
rect 120 93 122 107
rect 140 102 142 107
rect 145 105 147 107
rect 136 98 142 102
rect 140 93 142 98
rect 145 93 147 95
rect 163 93 165 107
rect 213 102 215 107
rect 218 102 220 104
rect 241 98 243 120
rect 213 96 215 98
rect 218 93 220 98
rect 241 92 243 94
rect 13 87 15 89
rect 29 85 31 89
rect 45 87 47 89
rect 68 87 70 89
rect 30 81 31 85
rect 73 84 75 89
rect 99 85 101 89
rect 120 87 122 89
rect 140 87 142 89
rect 29 78 31 81
rect 74 80 75 84
rect 100 81 101 85
rect 145 84 147 89
rect 163 87 165 89
rect 73 78 75 80
rect 99 77 101 81
rect 146 80 147 84
rect 145 78 147 80
rect 29 55 31 58
rect 73 56 75 58
rect 30 51 31 55
rect 74 52 75 56
rect 99 55 101 59
rect 145 56 147 58
rect 13 47 15 49
rect 29 47 31 51
rect 45 47 47 49
rect 68 47 70 49
rect 73 47 75 52
rect 100 51 101 55
rect 146 52 147 56
rect 290 55 292 58
rect 334 56 336 58
rect 99 47 101 51
rect 120 47 122 49
rect 140 47 142 49
rect 145 47 147 52
rect 291 51 292 55
rect 335 52 336 56
rect 360 55 362 59
rect 406 56 408 58
rect 163 47 165 49
rect 247 47 249 50
rect 265 47 267 50
rect 290 47 292 51
rect 306 47 308 49
rect 329 47 331 49
rect 334 47 336 52
rect 361 51 362 55
rect 407 52 408 56
rect 360 47 362 51
rect 381 47 383 49
rect 401 47 403 49
rect 406 47 408 52
rect 424 47 426 49
rect 13 29 15 43
rect 29 41 31 43
rect 29 29 31 31
rect 45 29 47 43
rect 68 38 70 43
rect 73 41 75 43
rect 99 41 101 43
rect 64 34 70 38
rect 68 29 70 34
rect 73 29 75 31
rect 99 29 101 31
rect 120 29 122 43
rect 140 38 142 43
rect 145 41 147 43
rect 136 34 142 38
rect 140 29 142 34
rect 145 29 147 31
rect 163 29 165 43
rect 213 40 215 43
rect 218 40 220 43
rect 247 38 249 43
rect 213 24 215 36
rect 218 34 220 36
rect 247 29 249 34
rect 265 29 267 43
rect 290 41 292 43
rect 290 29 292 31
rect 306 29 308 43
rect 329 38 331 43
rect 334 41 336 43
rect 360 41 362 43
rect 325 34 331 38
rect 329 29 331 34
rect 334 29 336 31
rect 360 29 362 31
rect 381 29 383 43
rect 401 38 403 43
rect 406 41 408 43
rect 397 34 403 38
rect 401 29 403 34
rect 406 29 408 31
rect 424 29 426 43
rect 218 24 220 26
rect 13 19 15 21
rect 29 18 31 21
rect 45 19 47 21
rect 68 19 70 21
rect 73 18 75 21
rect 99 18 101 21
rect 120 18 122 21
rect 140 19 142 21
rect 145 18 147 21
rect 163 19 165 21
rect 99 14 100 18
rect 247 18 249 21
rect 265 18 267 21
rect 290 18 292 21
rect 306 19 308 21
rect 329 19 331 21
rect 334 18 336 21
rect 360 18 362 21
rect 381 18 383 21
rect 401 19 403 21
rect 406 18 408 21
rect 424 19 426 21
rect 213 14 215 16
rect 29 11 31 14
rect 73 11 75 14
rect 99 11 101 14
rect 145 11 147 14
rect 218 11 220 16
rect 360 14 361 18
rect 290 11 292 14
rect 334 11 336 14
rect 360 11 362 14
rect 406 11 408 14
<< polycontact >>
rect 13 598 17 602
rect 50 598 54 602
rect 70 598 74 602
rect 108 598 112 602
rect 145 598 149 602
rect 182 598 186 602
rect 202 598 206 602
rect 240 598 244 602
rect 277 598 281 602
rect 314 598 318 602
rect 334 598 338 602
rect 372 598 376 602
rect 409 598 413 602
rect 446 598 450 602
rect 466 598 470 602
rect 504 598 508 602
rect 7 578 11 582
rect 25 580 29 584
rect 85 580 89 584
rect 43 571 47 578
rect 101 571 105 578
rect 122 575 126 579
rect 139 578 143 582
rect 157 580 161 584
rect 217 580 221 584
rect 175 571 179 578
rect 233 571 237 578
rect 254 575 258 579
rect 271 578 275 582
rect 289 580 293 584
rect 349 580 353 584
rect 307 571 311 578
rect 365 571 369 578
rect 386 575 390 579
rect 403 578 407 582
rect 421 580 425 584
rect 481 580 485 584
rect 439 571 443 578
rect 497 571 501 578
rect 518 575 522 579
rect 13 557 17 561
rect 50 555 54 559
rect 70 555 74 559
rect 106 555 110 559
rect 145 557 149 561
rect 182 555 186 559
rect 202 555 206 559
rect 238 555 242 559
rect 277 557 281 561
rect 314 555 318 559
rect 334 555 338 559
rect 370 555 374 559
rect 409 557 413 561
rect 446 555 450 559
rect 466 555 470 559
rect 502 555 506 559
rect 29 514 33 518
rect 73 514 77 518
rect 100 514 104 518
rect 145 514 149 518
rect 218 521 222 525
rect 183 507 187 511
rect 9 494 13 498
rect 41 495 45 499
rect 60 494 64 498
rect 116 495 120 499
rect 132 494 136 498
rect 159 494 163 498
rect 299 521 303 525
rect 210 503 214 507
rect 237 499 241 503
rect 264 507 268 511
rect 291 503 295 507
rect 318 499 322 503
rect 216 485 220 489
rect 297 485 301 489
rect 26 477 30 481
rect 70 476 74 480
rect 95 477 100 481
rect 142 476 146 480
rect 26 447 30 451
rect 70 448 74 452
rect 95 447 100 451
rect 142 448 146 452
rect 218 445 222 449
rect 299 445 303 449
rect 9 430 13 434
rect 41 429 45 433
rect 60 430 64 434
rect 116 429 120 433
rect 132 430 136 434
rect 159 430 163 434
rect 207 429 213 433
rect 288 429 294 433
rect 29 410 33 414
rect 73 410 77 414
rect 100 410 104 414
rect 145 410 149 414
rect 216 409 220 413
rect 297 409 301 413
rect 218 389 222 393
rect 29 382 33 386
rect 73 382 77 386
rect 100 382 104 386
rect 145 382 149 386
rect 323 389 327 393
rect 210 371 214 375
rect 9 362 13 366
rect 41 363 45 367
rect 60 362 64 366
rect 116 363 120 367
rect 132 362 136 366
rect 159 362 163 366
rect 237 367 241 371
rect 288 375 292 379
rect 315 371 319 375
rect 342 367 346 371
rect 216 353 220 357
rect 321 353 325 357
rect 26 345 30 349
rect 70 344 74 348
rect 95 345 100 349
rect 142 344 146 348
rect 26 315 30 319
rect 70 316 74 320
rect 95 315 100 319
rect 142 316 146 320
rect 218 314 222 318
rect 323 314 327 318
rect 9 298 13 302
rect 41 297 45 301
rect 60 298 64 302
rect 116 297 120 301
rect 132 298 136 302
rect 159 298 163 302
rect 207 298 213 302
rect 312 298 318 302
rect 29 278 33 282
rect 73 278 77 282
rect 100 278 104 282
rect 145 278 149 282
rect 216 278 220 282
rect 321 278 325 282
rect 218 257 222 261
rect 29 250 33 254
rect 73 250 77 254
rect 100 250 104 254
rect 145 250 149 254
rect 299 257 303 261
rect 210 239 214 243
rect 9 230 13 234
rect 41 231 45 235
rect 60 230 64 234
rect 116 231 120 235
rect 132 230 136 234
rect 159 230 163 234
rect 237 235 241 239
rect 264 243 268 247
rect 389 257 393 261
rect 291 239 295 243
rect 318 235 322 239
rect 354 243 358 247
rect 381 239 385 243
rect 408 235 412 239
rect 216 221 220 225
rect 297 221 301 225
rect 387 221 391 225
rect 26 213 30 217
rect 70 212 74 216
rect 95 213 100 217
rect 142 212 146 216
rect 26 183 30 187
rect 70 184 74 188
rect 95 183 100 187
rect 142 184 146 188
rect 218 179 222 183
rect 299 179 303 183
rect 389 179 393 183
rect 9 166 13 170
rect 41 165 45 169
rect 60 166 64 170
rect 116 165 120 169
rect 132 166 136 170
rect 159 166 163 170
rect 207 163 213 167
rect 288 163 294 167
rect 378 163 384 167
rect 29 146 33 150
rect 73 146 77 150
rect 100 146 104 150
rect 145 146 149 150
rect 216 143 220 147
rect 297 143 301 147
rect 387 143 391 147
rect 218 125 222 129
rect 29 118 33 122
rect 73 118 77 122
rect 100 118 104 122
rect 145 118 149 122
rect 210 107 214 111
rect 9 98 13 102
rect 41 99 45 103
rect 60 98 64 102
rect 116 99 120 103
rect 132 98 136 102
rect 159 98 163 102
rect 237 103 241 107
rect 216 89 220 93
rect 26 81 30 85
rect 70 80 74 84
rect 95 81 100 85
rect 142 80 146 84
rect 26 51 30 55
rect 70 52 74 56
rect 95 51 100 55
rect 142 52 146 56
rect 287 51 291 55
rect 331 52 335 56
rect 356 51 361 55
rect 403 52 407 56
rect 218 43 222 47
rect 9 34 13 38
rect 41 33 45 37
rect 60 34 64 38
rect 116 33 120 37
rect 132 34 136 38
rect 159 34 163 38
rect 207 27 213 31
rect 245 34 249 38
rect 302 33 306 37
rect 321 34 325 38
rect 377 33 381 37
rect 393 34 397 38
rect 420 34 424 38
rect 29 14 33 18
rect 73 14 77 18
rect 100 14 104 18
rect 145 14 149 18
rect 290 14 294 18
rect 334 14 338 18
rect 361 14 365 18
rect 406 14 410 18
rect 216 7 220 11
<< metal1 >>
rect -57 545 -53 623
rect -57 473 -53 541
rect -57 459 -53 469
rect -57 341 -53 455
rect -57 327 -53 337
rect -57 209 -53 323
rect -57 195 -53 205
rect -57 77 -53 191
rect -57 63 -53 73
rect -57 -21 -53 59
rect -57 -38 -53 -25
rect -43 616 -39 623
rect -43 612 9 616
rect 13 612 45 616
rect 49 612 112 616
rect 116 612 141 616
rect 145 612 177 616
rect 181 612 244 616
rect 248 612 273 616
rect 277 612 309 616
rect 313 612 376 616
rect 380 612 405 616
rect 409 612 441 616
rect 445 612 508 616
rect 512 612 528 616
rect -43 525 -39 612
rect 0 605 33 609
rect 37 605 61 609
rect 65 605 91 609
rect 95 605 128 609
rect 132 605 165 609
rect 169 605 193 609
rect 197 605 223 609
rect 227 605 260 609
rect 264 605 297 609
rect 301 605 325 609
rect 329 605 355 609
rect 359 605 392 609
rect 396 605 429 609
rect 433 605 457 609
rect 461 605 487 609
rect 491 605 524 609
rect 3 595 6 605
rect 24 595 27 605
rect 40 595 43 605
rect 54 598 59 602
rect 63 598 70 602
rect 82 595 85 605
rect 98 595 101 605
rect 119 595 122 605
rect 135 595 138 605
rect 156 595 159 605
rect 172 595 175 605
rect 186 598 191 602
rect 195 598 202 602
rect 214 595 217 605
rect 230 595 233 605
rect 251 595 254 605
rect 267 595 270 605
rect 288 595 291 605
rect 304 595 307 605
rect 318 598 323 602
rect 327 598 334 602
rect 346 595 349 605
rect 362 595 365 605
rect 383 595 386 605
rect 399 595 402 605
rect 420 595 423 605
rect 436 595 439 605
rect 450 598 455 602
rect 459 598 466 602
rect 478 595 481 605
rect 494 595 497 605
rect 515 595 518 605
rect 20 581 25 584
rect 29 581 53 584
rect 78 581 85 584
rect 89 581 111 584
rect 36 571 43 574
rect 47 575 66 578
rect 66 568 69 574
rect 94 571 101 574
rect 105 575 122 578
rect 152 581 157 584
rect 161 581 185 584
rect 210 581 217 584
rect 221 581 243 584
rect 168 571 175 574
rect 179 575 198 578
rect 198 568 201 574
rect 226 571 233 574
rect 237 575 254 578
rect 284 581 289 584
rect 293 581 317 584
rect 342 581 349 584
rect 353 581 375 584
rect 300 571 307 574
rect 311 575 330 578
rect 330 568 333 574
rect 358 571 365 574
rect 369 575 386 578
rect 416 581 421 584
rect 425 581 449 584
rect 474 581 481 584
rect 485 581 507 584
rect 432 571 439 574
rect 443 575 462 578
rect 3 552 6 564
rect 24 552 27 564
rect 40 552 43 564
rect 54 555 66 558
rect 82 552 85 564
rect 98 552 101 564
rect 119 552 122 564
rect 135 552 138 564
rect 156 552 159 564
rect 172 552 175 564
rect 186 555 198 558
rect 214 552 217 564
rect 230 552 233 564
rect 251 552 254 564
rect 267 552 270 564
rect 288 552 291 564
rect 304 552 307 564
rect 318 555 330 558
rect 346 552 349 564
rect 362 552 365 564
rect 383 552 386 564
rect 462 568 465 574
rect 490 571 497 574
rect 501 575 518 578
rect 399 552 402 564
rect 420 552 423 564
rect 436 552 439 564
rect 450 555 462 558
rect 478 552 481 564
rect 494 552 497 564
rect 515 552 518 564
rect 0 548 33 552
rect 37 548 61 552
rect 65 548 91 552
rect 95 548 165 552
rect 169 548 193 552
rect 197 548 223 552
rect 227 548 297 552
rect 301 548 325 552
rect 329 548 355 552
rect 359 548 429 552
rect 433 548 457 552
rect 461 548 487 552
rect 491 548 528 552
rect 0 541 9 545
rect 13 541 60 545
rect 64 541 110 545
rect 114 541 141 545
rect 145 541 192 545
rect 196 541 242 545
rect 246 541 273 545
rect 277 541 324 545
rect 328 541 374 545
rect 378 541 405 545
rect 409 541 456 545
rect 460 541 506 545
rect 510 541 528 545
rect 1 528 7 532
rect 11 528 23 532
rect 27 528 41 532
rect 45 528 52 532
rect 56 528 58 532
rect 62 528 77 532
rect 81 528 114 532
rect 118 528 119 532
rect 123 528 131 532
rect 135 528 159 532
rect 163 528 175 532
rect 179 528 199 532
rect 203 528 253 532
rect 257 528 280 532
rect 284 528 334 532
rect 338 528 357 532
rect -43 521 34 525
rect 38 521 65 525
rect 69 521 87 525
rect 91 521 152 525
rect 156 521 170 525
rect 182 524 185 528
rect -43 407 -39 521
rect 77 514 80 518
rect 104 514 105 518
rect 149 514 151 518
rect 191 511 194 516
rect 206 518 209 528
rect 236 524 239 528
rect 263 524 266 528
rect 6 494 9 497
rect 17 497 20 503
rect 24 497 27 503
rect 17 494 27 497
rect 17 489 20 494
rect 24 489 27 494
rect 33 499 36 503
rect 33 495 35 499
rect 39 495 41 499
rect 49 498 52 503
rect 77 500 80 503
rect 49 496 60 498
rect 33 489 36 495
rect 49 494 55 496
rect 49 489 52 494
rect 59 494 60 496
rect 78 496 80 500
rect 77 489 80 496
rect 180 507 183 510
rect 222 507 225 510
rect 93 499 96 503
rect 103 499 106 503
rect 103 495 112 499
rect 124 498 127 503
rect 149 499 152 503
rect 93 489 96 495
rect 103 489 106 495
rect 124 494 125 498
rect 129 494 132 497
rect 151 495 152 499
rect 167 498 170 503
rect 191 502 194 507
rect 199 503 210 506
rect 222 504 230 507
rect 124 489 127 494
rect 149 489 152 495
rect 167 489 170 494
rect 69 476 70 480
rect 94 477 95 481
rect 141 476 142 480
rect 1 469 22 473
rect 26 469 81 473
rect 85 469 106 473
rect 110 469 137 473
rect 141 469 170 473
rect 182 466 185 498
rect 199 497 202 503
rect 222 498 225 504
rect 234 499 237 502
rect 245 502 248 516
rect 272 511 275 516
rect 287 518 290 528
rect 317 524 320 528
rect 256 507 257 510
rect 261 507 264 510
rect 303 507 306 510
rect 245 499 253 502
rect 272 502 275 507
rect 245 494 248 499
rect 253 495 257 499
rect 280 503 291 506
rect 303 504 311 507
rect 197 488 202 493
rect 206 466 209 494
rect 236 466 239 490
rect 263 466 266 498
rect 280 497 283 503
rect 303 498 306 504
rect 315 499 318 502
rect 326 502 329 516
rect 326 499 338 502
rect 326 494 329 499
rect 278 488 283 493
rect 287 466 290 494
rect 317 466 320 490
rect 1 462 8 466
rect 12 462 14 466
rect 18 462 22 466
rect 26 462 40 466
rect 44 462 49 466
rect 53 462 58 466
rect 62 462 81 466
rect 85 462 115 466
rect 119 462 130 466
rect 134 462 158 466
rect 162 462 175 466
rect 179 462 199 466
rect 203 462 253 466
rect 260 462 280 466
rect 284 462 334 466
rect 1 455 22 459
rect 26 455 81 459
rect 85 455 106 459
rect 110 455 137 459
rect 141 455 170 459
rect 69 448 70 452
rect 94 447 95 451
rect 141 448 142 452
rect 17 434 20 439
rect 24 434 27 439
rect 7 431 9 434
rect 17 431 27 434
rect 17 425 20 431
rect 24 425 27 431
rect 33 433 36 439
rect 49 434 52 439
rect 33 429 35 433
rect 39 429 41 433
rect 49 432 55 434
rect 59 432 60 434
rect 49 430 60 432
rect 77 432 80 439
rect 33 425 36 429
rect 49 425 52 430
rect 78 428 80 432
rect 77 425 80 428
rect 93 433 96 439
rect 103 433 106 439
rect 124 434 127 439
rect 103 429 112 433
rect 124 430 125 434
rect 129 431 132 434
rect 149 433 152 439
rect 167 434 170 439
rect 206 442 209 462
rect 287 442 290 462
rect 93 425 96 429
rect 103 425 106 429
rect 124 425 127 430
rect 151 429 152 433
rect 149 425 152 429
rect 167 425 170 430
rect 197 429 202 434
rect 206 430 207 433
rect 222 432 225 438
rect 222 429 230 432
rect 277 429 282 434
rect 286 430 288 433
rect 303 432 306 438
rect 303 429 311 432
rect 222 426 225 429
rect 303 426 306 429
rect 77 410 80 414
rect 104 410 105 414
rect 149 410 151 414
rect -43 403 34 407
rect 38 403 65 407
rect 69 403 87 407
rect 91 403 152 407
rect 156 403 170 407
rect -43 393 -39 403
rect 206 400 209 418
rect 287 400 290 418
rect 1 396 7 400
rect 11 396 23 400
rect 27 396 41 400
rect 45 396 52 400
rect 56 396 58 400
rect 62 396 77 400
rect 81 396 114 400
rect 118 396 119 400
rect 123 396 131 400
rect 135 396 159 400
rect 163 396 175 400
rect 179 396 199 400
rect 203 396 253 400
rect 257 396 280 400
rect 284 396 342 400
rect 346 396 357 400
rect -43 389 34 393
rect 38 389 65 393
rect 69 389 87 393
rect 91 389 152 393
rect 156 389 170 393
rect -43 275 -39 389
rect 206 386 209 396
rect 236 392 239 396
rect 287 392 290 396
rect 77 382 80 386
rect 104 382 105 386
rect 149 382 151 386
rect 6 362 9 365
rect 17 365 20 371
rect 24 365 27 371
rect 17 362 27 365
rect 17 357 20 362
rect 24 357 27 362
rect 33 367 36 371
rect 33 363 35 367
rect 39 363 41 367
rect 49 366 52 371
rect 77 368 80 371
rect 49 364 60 366
rect 33 357 36 363
rect 49 362 55 364
rect 49 357 52 362
rect 59 362 60 364
rect 78 364 80 368
rect 77 357 80 364
rect 222 375 225 378
rect 93 367 96 371
rect 103 367 106 371
rect 103 363 112 367
rect 124 366 127 371
rect 149 367 152 371
rect 93 357 96 363
rect 103 357 106 363
rect 124 362 125 366
rect 129 362 132 365
rect 151 363 152 367
rect 167 366 170 371
rect 199 371 210 374
rect 222 372 230 375
rect 124 357 127 362
rect 149 357 152 363
rect 199 365 202 371
rect 222 366 225 372
rect 234 367 237 370
rect 245 370 248 384
rect 296 379 299 384
rect 311 386 314 396
rect 341 392 344 396
rect 280 375 281 378
rect 285 375 288 378
rect 327 375 330 378
rect 253 370 258 375
rect 296 370 299 375
rect 245 367 253 370
rect 167 357 170 362
rect 245 362 248 367
rect 304 371 315 374
rect 327 372 335 375
rect 197 356 202 361
rect 69 344 70 348
rect 94 345 95 349
rect 141 344 142 348
rect 1 337 22 341
rect 26 337 81 341
rect 85 337 106 341
rect 110 337 137 341
rect 141 337 170 341
rect 206 334 209 362
rect 236 334 239 358
rect 287 334 290 366
rect 304 365 307 371
rect 327 366 330 372
rect 339 367 342 370
rect 350 370 353 384
rect 350 367 356 370
rect 350 362 353 367
rect 302 356 307 361
rect 311 334 314 362
rect 341 334 344 358
rect 1 330 8 334
rect 12 330 14 334
rect 18 330 22 334
rect 26 330 40 334
rect 44 330 49 334
rect 53 330 58 334
rect 62 330 81 334
rect 85 330 115 334
rect 119 330 130 334
rect 134 330 158 334
rect 162 330 175 334
rect 179 330 199 334
rect 203 330 253 334
rect 257 330 280 334
rect 284 330 304 334
rect 308 330 356 334
rect 1 323 22 327
rect 26 323 81 327
rect 85 323 106 327
rect 110 323 137 327
rect 141 323 170 327
rect 69 316 70 320
rect 94 315 95 319
rect 141 316 142 320
rect 206 311 209 330
rect 311 311 314 330
rect 17 302 20 307
rect 24 302 27 307
rect 7 299 9 302
rect 17 299 27 302
rect 17 293 20 299
rect 24 293 27 299
rect 33 301 36 307
rect 49 302 52 307
rect 33 297 35 301
rect 39 297 41 301
rect 49 300 55 302
rect 59 300 60 302
rect 49 298 60 300
rect 77 300 80 307
rect 33 293 36 297
rect 49 293 52 298
rect 78 296 80 300
rect 77 293 80 296
rect 93 301 96 307
rect 103 301 106 307
rect 124 302 127 307
rect 103 297 112 301
rect 124 298 125 302
rect 129 299 132 302
rect 149 301 152 307
rect 167 302 170 307
rect 93 293 96 297
rect 103 293 106 297
rect 124 293 127 298
rect 151 297 152 301
rect 196 298 201 303
rect 205 299 207 302
rect 222 301 225 307
rect 222 298 230 301
rect 302 298 307 303
rect 311 299 312 302
rect 327 301 330 307
rect 327 298 335 301
rect 149 293 152 297
rect 167 293 170 298
rect 222 295 225 298
rect 327 295 330 298
rect 77 278 80 282
rect 104 278 105 282
rect 149 278 151 282
rect -43 271 34 275
rect 38 271 65 275
rect 69 271 87 275
rect 91 271 152 275
rect 156 271 170 275
rect -43 261 -39 271
rect 206 268 209 287
rect 311 268 314 287
rect 1 264 7 268
rect 11 264 23 268
rect 27 264 41 268
rect 45 264 52 268
rect 56 264 58 268
rect 62 264 77 268
rect 81 264 114 268
rect 118 264 119 268
rect 123 264 131 268
rect 135 264 159 268
rect 163 264 175 268
rect 179 264 199 268
rect 203 264 253 268
rect 257 264 280 268
rect 284 264 334 268
rect 338 264 342 268
rect 346 264 370 268
rect 374 264 424 268
rect -43 257 34 261
rect 38 257 65 261
rect 69 257 87 261
rect 91 257 152 261
rect 156 257 170 261
rect -43 143 -39 257
rect 206 254 209 264
rect 236 260 239 264
rect 263 260 266 264
rect 77 250 80 254
rect 104 250 105 254
rect 149 250 151 254
rect 6 230 9 233
rect 17 233 20 239
rect 24 233 27 239
rect 17 230 27 233
rect 17 225 20 230
rect 24 225 27 230
rect 33 235 36 239
rect 33 231 35 235
rect 39 231 41 235
rect 49 234 52 239
rect 77 236 80 239
rect 49 232 60 234
rect 33 225 36 231
rect 49 230 55 232
rect 49 225 52 230
rect 59 230 60 232
rect 78 232 80 236
rect 77 225 80 232
rect 222 243 225 246
rect 93 235 96 239
rect 103 235 106 239
rect 103 231 112 235
rect 124 234 127 239
rect 149 235 152 239
rect 93 225 96 231
rect 103 225 106 231
rect 124 230 125 234
rect 129 230 132 233
rect 151 231 152 235
rect 167 234 170 239
rect 199 239 210 242
rect 222 240 230 243
rect 124 225 127 230
rect 149 225 152 231
rect 199 233 202 239
rect 222 234 225 240
rect 234 235 237 238
rect 245 238 248 252
rect 272 247 275 252
rect 287 254 290 264
rect 317 260 320 264
rect 353 260 356 264
rect 256 243 257 246
rect 261 243 264 246
rect 303 243 306 246
rect 245 235 253 238
rect 272 238 275 243
rect 167 225 170 230
rect 245 230 248 235
rect 253 231 257 235
rect 280 239 291 242
rect 303 240 311 243
rect 197 224 202 229
rect 69 212 70 216
rect 94 213 95 217
rect 141 212 142 216
rect 1 205 22 209
rect 26 205 81 209
rect 85 205 106 209
rect 110 205 137 209
rect 141 205 170 209
rect 206 202 209 230
rect 236 202 239 226
rect 263 202 266 234
rect 280 233 283 239
rect 303 234 306 240
rect 315 235 318 238
rect 326 238 329 252
rect 362 247 365 252
rect 377 254 380 264
rect 407 260 410 264
rect 351 243 354 246
rect 393 243 396 246
rect 326 235 335 238
rect 362 238 365 243
rect 326 230 329 235
rect 278 224 283 229
rect 287 202 290 230
rect 369 241 381 242
rect 373 239 381 241
rect 393 240 401 243
rect 393 234 396 240
rect 405 235 408 238
rect 416 238 419 252
rect 416 235 428 238
rect 317 202 320 226
rect 353 202 356 234
rect 416 230 419 235
rect 377 202 380 230
rect 407 202 410 226
rect 1 198 8 202
rect 12 198 14 202
rect 18 198 22 202
rect 26 198 40 202
rect 44 198 49 202
rect 53 198 58 202
rect 62 198 81 202
rect 85 198 115 202
rect 119 198 130 202
rect 134 198 158 202
rect 162 198 175 202
rect 179 198 199 202
rect 203 198 253 202
rect 260 198 280 202
rect 284 198 334 202
rect 338 198 370 202
rect 374 198 424 202
rect 1 191 22 195
rect 26 191 81 195
rect 85 191 106 195
rect 110 191 137 195
rect 141 191 170 195
rect 69 184 70 188
rect 94 183 95 187
rect 141 184 142 188
rect 17 170 20 175
rect 24 170 27 175
rect 7 167 9 170
rect 17 167 27 170
rect 17 161 20 167
rect 24 161 27 167
rect 33 169 36 175
rect 49 170 52 175
rect 33 165 35 169
rect 39 165 41 169
rect 49 168 55 170
rect 59 168 60 170
rect 49 166 60 168
rect 77 168 80 175
rect 33 161 36 165
rect 49 161 52 166
rect 78 164 80 168
rect 77 161 80 164
rect 93 169 96 175
rect 103 169 106 175
rect 124 170 127 175
rect 103 165 112 169
rect 124 166 125 170
rect 129 167 132 170
rect 149 169 152 175
rect 167 170 170 175
rect 206 176 209 198
rect 287 176 290 198
rect 377 176 380 198
rect 93 161 96 165
rect 103 161 106 165
rect 124 161 127 166
rect 151 165 152 169
rect 149 161 152 165
rect 167 161 170 166
rect 197 163 202 168
rect 206 164 207 167
rect 222 166 225 172
rect 222 163 230 166
rect 277 163 282 168
rect 286 164 288 167
rect 303 166 306 172
rect 303 163 311 166
rect 370 164 378 167
rect 393 166 396 172
rect 393 163 401 166
rect 222 160 225 163
rect 303 160 306 163
rect 393 160 396 163
rect 77 146 80 150
rect 104 146 105 150
rect 149 146 151 150
rect -43 139 34 143
rect 38 139 65 143
rect 69 139 87 143
rect 91 139 152 143
rect 156 139 170 143
rect -43 129 -39 139
rect 206 136 209 152
rect 287 136 290 152
rect 377 136 380 152
rect 1 132 7 136
rect 11 132 23 136
rect 27 132 41 136
rect 45 132 52 136
rect 56 132 58 136
rect 62 132 77 136
rect 81 132 114 136
rect 118 132 119 136
rect 123 132 131 136
rect 135 132 159 136
rect 163 132 175 136
rect 179 132 199 136
rect 203 132 253 136
rect 257 132 280 136
rect 284 132 370 136
rect 374 132 428 136
rect -43 125 34 129
rect 38 125 65 129
rect 69 125 87 129
rect 91 125 152 129
rect 156 125 170 129
rect -43 11 -39 125
rect 206 122 209 132
rect 236 128 239 132
rect 77 118 80 122
rect 104 118 105 122
rect 149 118 151 122
rect 6 98 9 101
rect 17 101 20 107
rect 24 101 27 107
rect 17 98 27 101
rect 17 93 20 98
rect 24 93 27 98
rect 33 103 36 107
rect 33 99 35 103
rect 39 99 41 103
rect 49 102 52 107
rect 77 104 80 107
rect 49 100 60 102
rect 33 93 36 99
rect 49 98 55 100
rect 49 93 52 98
rect 59 98 60 100
rect 78 100 80 104
rect 77 93 80 100
rect 222 111 225 114
rect 93 103 96 107
rect 103 103 106 107
rect 103 99 112 103
rect 124 102 127 107
rect 149 103 152 107
rect 93 93 96 99
rect 103 93 106 99
rect 124 98 125 102
rect 129 98 132 101
rect 151 99 152 103
rect 167 102 170 107
rect 199 107 210 110
rect 222 108 230 111
rect 124 93 127 98
rect 149 93 152 99
rect 199 101 202 107
rect 222 102 225 108
rect 234 103 237 106
rect 245 106 248 120
rect 253 106 258 111
rect 245 103 253 106
rect 167 93 170 98
rect 245 98 248 103
rect 197 92 202 97
rect 69 80 70 84
rect 94 81 95 85
rect 141 80 142 84
rect 1 73 22 77
rect 26 73 81 77
rect 85 73 106 77
rect 110 73 137 77
rect 141 73 170 77
rect 206 70 209 98
rect 236 70 239 94
rect 1 66 8 70
rect 12 66 14 70
rect 18 66 22 70
rect 26 66 40 70
rect 44 66 49 70
rect 53 66 58 70
rect 62 66 81 70
rect 85 66 115 70
rect 119 66 130 70
rect 134 66 158 70
rect 162 66 175 70
rect 179 66 199 70
rect 203 66 283 70
rect 287 66 301 70
rect 305 66 310 70
rect 314 66 319 70
rect 323 66 342 70
rect 346 66 376 70
rect 380 66 391 70
rect 395 66 419 70
rect 423 66 432 70
rect 1 59 22 63
rect 26 59 81 63
rect 85 59 106 63
rect 110 59 137 63
rect 141 59 170 63
rect 69 52 70 56
rect 94 51 95 55
rect 141 52 142 56
rect 17 38 20 43
rect 24 38 27 43
rect 7 35 9 38
rect 17 35 27 38
rect 17 29 20 35
rect 24 29 27 35
rect 33 37 36 43
rect 49 38 52 43
rect 33 33 35 37
rect 39 33 41 37
rect 49 36 55 38
rect 59 36 60 38
rect 49 34 60 36
rect 77 36 80 43
rect 33 29 36 33
rect 49 29 52 34
rect 78 32 80 36
rect 77 29 80 32
rect 93 37 96 43
rect 103 37 106 43
rect 124 38 127 43
rect 103 33 112 37
rect 124 34 125 38
rect 129 35 132 38
rect 149 37 152 43
rect 167 38 170 43
rect 206 40 209 66
rect 242 59 261 63
rect 265 59 283 63
rect 287 59 342 63
rect 346 59 367 63
rect 371 59 398 63
rect 402 59 431 63
rect 242 47 245 59
rect 330 52 331 56
rect 355 51 356 55
rect 402 52 403 56
rect 93 29 96 33
rect 103 29 106 33
rect 124 29 127 34
rect 151 33 152 37
rect 269 38 272 43
rect 278 38 281 43
rect 285 38 288 43
rect 149 29 152 33
rect 167 29 170 34
rect 196 27 201 32
rect 205 28 207 31
rect 222 30 225 36
rect 254 35 288 38
rect 222 27 230 30
rect 222 24 225 27
rect 77 14 80 18
rect 104 14 105 18
rect 149 14 151 18
rect 254 21 257 35
rect 278 29 281 35
rect 285 29 288 35
rect 294 37 297 43
rect 310 38 313 43
rect 294 33 296 37
rect 300 33 302 37
rect 310 36 316 38
rect 320 36 321 38
rect 310 34 321 36
rect 338 36 341 43
rect 294 29 297 33
rect 310 29 313 34
rect 339 32 341 36
rect 338 29 341 32
rect 354 37 357 43
rect 364 37 367 43
rect 385 38 388 43
rect 364 33 373 37
rect 385 34 386 38
rect 390 35 393 38
rect 410 37 413 43
rect 428 38 431 43
rect 354 29 357 33
rect 364 29 367 33
rect 385 29 388 34
rect 412 33 413 37
rect 410 29 413 33
rect 428 29 431 34
rect -43 7 34 11
rect 38 7 65 11
rect 69 7 87 11
rect 91 7 152 11
rect 156 7 170 11
rect -43 -14 -39 7
rect 206 4 209 16
rect 338 14 341 18
rect 365 14 366 18
rect 410 14 412 18
rect 246 7 251 11
rect 255 7 295 11
rect 299 7 326 11
rect 330 7 348 11
rect 352 7 413 11
rect 417 7 431 11
rect 1 0 7 4
rect 11 0 23 4
rect 27 0 41 4
rect 45 0 52 4
rect 56 0 58 4
rect 62 0 77 4
rect 81 0 114 4
rect 118 0 119 4
rect 123 0 131 4
rect 135 0 159 4
rect 163 0 199 4
rect 203 0 242 4
rect 246 0 253 4
rect 257 0 268 4
rect 272 0 284 4
rect 288 0 302 4
rect 306 0 313 4
rect 317 0 319 4
rect 323 0 338 4
rect 342 0 375 4
rect 379 0 380 4
rect 384 0 392 4
rect 396 0 420 4
rect 424 0 432 4
rect -43 -17 250 -14
rect -43 -38 -39 -17
rect -26 -24 260 -21
<< m2contact >>
rect -57 541 -53 545
rect -57 469 -53 473
rect -57 455 -53 459
rect -57 337 -53 341
rect -57 323 -53 327
rect -57 205 -53 209
rect -57 191 -53 195
rect -57 73 -53 77
rect -57 59 -53 63
rect -57 -25 -53 -21
rect 9 612 13 616
rect 45 612 49 616
rect 112 612 116 616
rect 141 612 145 616
rect 177 612 181 616
rect 244 612 248 616
rect 273 612 277 616
rect 309 612 313 616
rect 376 612 380 616
rect 405 612 409 616
rect 441 612 445 616
rect 508 612 512 616
rect 9 598 13 602
rect 59 598 63 602
rect 112 598 116 602
rect 141 598 145 602
rect 191 598 195 602
rect 244 598 248 602
rect 273 598 277 602
rect 323 598 327 602
rect 376 598 380 602
rect 405 598 409 602
rect 455 598 459 602
rect 508 598 512 602
rect 32 587 36 591
rect 3 578 7 582
rect 16 581 20 587
rect 53 581 57 587
rect 66 583 70 587
rect 90 587 94 591
rect 164 587 168 591
rect 74 581 78 587
rect 111 581 115 587
rect 127 583 131 587
rect 16 568 20 572
rect 32 568 36 574
rect 66 574 70 578
rect 53 568 57 572
rect 74 568 78 572
rect 90 568 94 574
rect 135 578 139 582
rect 148 581 152 587
rect 185 581 189 587
rect 198 583 202 587
rect 222 587 226 591
rect 296 587 300 591
rect 206 581 210 587
rect 243 581 247 587
rect 259 583 263 587
rect 111 568 115 572
rect 127 568 131 572
rect 148 568 152 572
rect 164 568 168 574
rect 198 574 202 578
rect 185 568 189 572
rect 206 568 210 572
rect 222 568 226 574
rect 267 578 271 582
rect 280 581 284 587
rect 317 581 321 587
rect 330 583 334 587
rect 354 587 358 591
rect 428 587 432 591
rect 338 581 342 587
rect 375 581 379 587
rect 391 583 395 587
rect 243 568 247 572
rect 259 568 263 572
rect 280 568 284 572
rect 296 568 300 574
rect 330 574 334 578
rect 317 568 321 572
rect 338 568 342 572
rect 354 568 358 574
rect 399 578 403 582
rect 412 581 416 587
rect 449 581 453 587
rect 462 583 466 587
rect 486 587 490 591
rect 470 581 474 587
rect 507 581 511 587
rect 523 583 527 587
rect 375 568 379 572
rect 391 568 395 572
rect 412 568 416 572
rect 428 568 432 574
rect 462 574 466 578
rect 449 568 453 572
rect 9 557 13 561
rect 46 555 50 559
rect 66 555 70 559
rect 110 555 114 559
rect 141 557 145 561
rect 178 555 182 559
rect 198 555 202 559
rect 242 555 246 559
rect 273 557 277 561
rect 310 555 314 559
rect 330 555 334 559
rect 374 555 378 559
rect 391 560 395 564
rect 470 568 474 572
rect 486 568 490 574
rect 507 568 511 572
rect 523 568 527 572
rect 405 557 409 561
rect 442 555 446 559
rect 462 555 466 559
rect 506 555 510 559
rect 523 560 527 564
rect -4 541 0 545
rect 9 541 13 545
rect 60 541 64 545
rect 110 541 114 545
rect 141 541 145 545
rect 192 541 196 545
rect 242 541 246 545
rect 273 541 277 545
rect 324 541 328 545
rect 374 541 378 545
rect 405 541 409 545
rect 456 541 460 545
rect 506 541 510 545
rect 7 528 11 532
rect 41 528 45 532
rect 58 528 62 532
rect 114 528 118 532
rect 131 528 135 532
rect 159 528 163 532
rect 34 521 38 525
rect 65 521 69 525
rect 87 521 91 525
rect 152 521 156 525
rect 8 511 12 515
rect 33 514 37 518
rect 40 511 44 515
rect 58 511 62 515
rect 80 514 84 518
rect 105 514 109 518
rect 115 511 119 515
rect 131 511 135 515
rect 151 514 155 518
rect 158 511 162 515
rect 222 521 226 525
rect 2 494 6 498
rect 35 495 39 499
rect 55 492 59 496
rect 74 496 78 500
rect 176 507 180 511
rect 191 507 195 511
rect 93 495 97 499
rect 112 495 116 499
rect 125 494 129 498
rect 147 495 151 499
rect 155 494 159 498
rect 167 494 171 498
rect 8 481 12 485
rect 40 481 44 485
rect 58 481 62 485
rect 115 481 119 485
rect 130 481 134 485
rect 158 481 162 485
rect 22 477 26 481
rect 65 476 69 480
rect 87 477 94 481
rect 137 476 141 480
rect -3 469 1 473
rect 22 469 26 473
rect 81 469 85 473
rect 106 469 110 473
rect 137 469 141 473
rect 230 499 234 507
rect 303 521 307 525
rect 257 507 261 511
rect 272 507 276 511
rect 253 499 257 503
rect 199 493 203 497
rect 212 485 216 489
rect 311 499 315 507
rect 338 499 342 503
rect 280 493 284 497
rect 293 485 297 489
rect 8 462 12 466
rect 22 462 26 466
rect 40 462 44 466
rect 58 462 62 466
rect 81 462 85 466
rect 115 462 119 466
rect 130 462 134 466
rect 158 462 162 466
rect -3 455 1 459
rect 22 455 26 459
rect 81 455 85 459
rect 106 455 110 459
rect 137 455 141 459
rect 22 447 26 451
rect 65 448 69 452
rect 87 447 94 451
rect 137 448 141 452
rect 8 443 12 447
rect 40 443 44 447
rect 58 443 62 447
rect 115 443 119 447
rect 130 443 134 447
rect 158 443 162 447
rect 3 431 7 435
rect 35 429 39 433
rect 55 432 59 436
rect 74 428 78 432
rect 93 429 97 433
rect 112 429 116 433
rect 125 430 129 434
rect 222 445 226 449
rect 303 445 307 449
rect 147 429 151 433
rect 155 430 159 434
rect 167 430 171 434
rect 202 430 206 434
rect 230 429 234 433
rect 282 430 286 434
rect 311 429 315 433
rect 8 413 12 417
rect 33 410 37 414
rect 40 413 44 417
rect 58 413 62 417
rect 80 410 84 414
rect 105 410 109 414
rect 115 413 119 417
rect 131 413 135 417
rect 151 410 155 414
rect 158 413 162 417
rect 34 403 38 407
rect 65 403 69 407
rect 87 403 91 407
rect 152 403 156 407
rect 212 409 216 413
rect 293 409 297 413
rect 7 396 11 400
rect 41 396 45 400
rect 58 396 62 400
rect 114 396 118 400
rect 131 396 135 400
rect 159 396 163 400
rect 34 389 38 393
rect 65 389 69 393
rect 87 389 91 393
rect 152 389 156 393
rect 222 389 226 393
rect 8 379 12 383
rect 33 382 37 386
rect 40 379 44 383
rect 58 379 62 383
rect 80 382 84 386
rect 105 382 109 386
rect 115 379 119 383
rect 131 379 135 383
rect 151 382 155 386
rect 158 379 162 383
rect 2 362 6 366
rect 35 363 39 367
rect 55 360 59 364
rect 74 364 78 368
rect 93 363 97 367
rect 112 363 116 367
rect 125 362 129 366
rect 147 363 151 367
rect 155 362 159 366
rect 167 362 171 366
rect 230 367 234 375
rect 327 389 331 393
rect 281 375 285 379
rect 296 375 300 379
rect 199 361 203 365
rect 253 366 257 370
rect 8 349 12 353
rect 40 349 44 353
rect 58 349 62 353
rect 115 349 119 353
rect 130 349 134 353
rect 158 349 162 353
rect 22 345 26 349
rect 65 344 69 348
rect 87 345 94 349
rect 137 344 141 348
rect -3 337 1 341
rect 22 337 26 341
rect 81 337 85 341
rect 106 337 110 341
rect 137 337 141 341
rect 212 353 216 357
rect 335 367 339 375
rect 356 367 360 371
rect 304 361 308 365
rect 317 353 321 357
rect 8 330 12 334
rect 22 330 26 334
rect 40 330 44 334
rect 58 330 62 334
rect 81 330 85 334
rect 115 330 119 334
rect 130 330 134 334
rect 158 330 162 334
rect -3 323 1 327
rect 22 323 26 327
rect 81 323 85 327
rect 106 323 110 327
rect 137 323 141 327
rect 22 315 26 319
rect 65 316 69 320
rect 87 315 94 319
rect 137 316 141 320
rect 8 311 12 315
rect 40 311 44 315
rect 58 311 62 315
rect 115 311 119 315
rect 130 311 134 315
rect 158 311 162 315
rect 222 314 226 318
rect 327 314 331 318
rect 3 299 7 303
rect 35 297 39 301
rect 55 300 59 304
rect 74 296 78 300
rect 93 297 97 301
rect 112 297 116 301
rect 125 298 129 302
rect 147 297 151 301
rect 155 298 159 302
rect 167 298 171 302
rect 201 299 205 303
rect 230 298 234 302
rect 307 299 311 303
rect 335 298 339 302
rect 8 281 12 285
rect 33 278 37 282
rect 40 281 44 285
rect 58 281 62 285
rect 80 278 84 282
rect 105 278 109 282
rect 115 281 119 285
rect 131 281 135 285
rect 151 278 155 282
rect 158 281 162 285
rect 34 271 38 275
rect 65 271 69 275
rect 87 271 91 275
rect 152 271 156 275
rect 212 278 216 282
rect 317 278 321 282
rect 7 264 11 268
rect 41 264 45 268
rect 58 264 62 268
rect 114 264 118 268
rect 131 264 135 268
rect 159 264 163 268
rect 34 257 38 261
rect 65 257 69 261
rect 87 257 91 261
rect 152 257 156 261
rect 222 257 226 261
rect 8 247 12 251
rect 33 250 37 254
rect 40 247 44 251
rect 58 247 62 251
rect 80 250 84 254
rect 105 250 109 254
rect 115 247 119 251
rect 131 247 135 251
rect 151 250 155 254
rect 158 247 162 251
rect 2 230 6 234
rect 35 231 39 235
rect 55 228 59 232
rect 74 232 78 236
rect 93 231 97 235
rect 112 231 116 235
rect 125 230 129 234
rect 147 231 151 235
rect 155 230 159 234
rect 167 230 171 234
rect 230 235 234 243
rect 303 257 307 261
rect 257 243 261 247
rect 272 243 276 247
rect 253 235 257 239
rect 199 229 203 233
rect 8 217 12 221
rect 40 217 44 221
rect 58 217 62 221
rect 115 217 119 221
rect 130 217 134 221
rect 158 217 162 221
rect 22 213 26 217
rect 65 212 69 216
rect 87 213 94 217
rect 137 212 141 216
rect -3 205 1 209
rect 22 205 26 209
rect 81 205 85 209
rect 106 205 110 209
rect 137 205 141 209
rect 212 221 216 225
rect 311 235 315 243
rect 393 257 397 261
rect 347 243 351 247
rect 362 243 366 247
rect 335 235 339 239
rect 280 229 284 233
rect 369 237 373 241
rect 401 235 405 243
rect 425 238 429 242
rect 293 221 297 225
rect 383 221 387 225
rect 8 198 12 202
rect 22 198 26 202
rect 40 198 44 202
rect 58 198 62 202
rect 81 198 85 202
rect 115 198 119 202
rect 130 198 134 202
rect 158 198 162 202
rect -3 191 1 195
rect 22 191 26 195
rect 81 191 85 195
rect 106 191 110 195
rect 137 191 141 195
rect 22 183 26 187
rect 65 184 69 188
rect 87 183 94 187
rect 137 184 141 188
rect 8 179 12 183
rect 40 179 44 183
rect 58 179 62 183
rect 115 179 119 183
rect 130 179 134 183
rect 158 179 162 183
rect 3 167 7 171
rect 35 165 39 169
rect 55 168 59 172
rect 74 164 78 168
rect 93 165 97 169
rect 112 165 116 169
rect 125 166 129 170
rect 222 179 226 183
rect 303 179 307 183
rect 393 179 397 183
rect 147 165 151 169
rect 155 166 159 170
rect 167 166 171 170
rect 202 164 206 168
rect 230 163 234 167
rect 282 164 286 168
rect 311 163 315 167
rect 366 164 370 168
rect 401 163 405 167
rect 8 149 12 153
rect 33 146 37 150
rect 40 149 44 153
rect 58 149 62 153
rect 80 146 84 150
rect 105 146 109 150
rect 115 149 119 153
rect 131 149 135 153
rect 151 146 155 150
rect 158 149 162 153
rect 34 139 38 143
rect 65 139 69 143
rect 87 139 91 143
rect 152 139 156 143
rect 212 143 216 147
rect 293 143 297 147
rect 383 143 387 147
rect 7 132 11 136
rect 41 132 45 136
rect 58 132 62 136
rect 114 132 118 136
rect 131 132 135 136
rect 159 132 163 136
rect 34 125 38 129
rect 65 125 69 129
rect 87 125 91 129
rect 152 125 156 129
rect 222 125 226 129
rect 8 115 12 119
rect 33 118 37 122
rect 40 115 44 119
rect 58 115 62 119
rect 80 118 84 122
rect 105 118 109 122
rect 115 115 119 119
rect 131 115 135 119
rect 151 118 155 122
rect 158 115 162 119
rect 2 98 6 102
rect 35 99 39 103
rect 55 96 59 100
rect 74 100 78 104
rect 93 99 97 103
rect 112 99 116 103
rect 125 98 129 102
rect 147 99 151 103
rect 155 98 159 102
rect 167 98 171 102
rect 230 103 234 111
rect 199 97 203 101
rect 253 102 257 106
rect 8 85 12 89
rect 40 85 44 89
rect 58 85 62 89
rect 115 85 119 89
rect 130 85 134 89
rect 158 85 162 89
rect 22 81 26 85
rect 65 80 69 84
rect 87 81 94 85
rect 137 80 141 84
rect -3 73 1 77
rect 22 73 26 77
rect 81 73 85 77
rect 106 73 110 77
rect 137 73 141 77
rect 212 89 216 93
rect 8 66 12 70
rect 22 66 26 70
rect 40 66 44 70
rect 58 66 62 70
rect 81 66 85 70
rect 115 66 119 70
rect 130 66 134 70
rect 158 66 162 70
rect 283 66 287 70
rect 301 66 305 70
rect 319 66 323 70
rect 342 66 346 70
rect 376 66 380 70
rect 391 66 395 70
rect 419 66 423 70
rect -3 59 1 63
rect 22 59 26 63
rect 81 59 85 63
rect 106 59 110 63
rect 137 59 141 63
rect 22 51 26 55
rect 65 52 69 56
rect 87 51 94 55
rect 137 52 141 56
rect 8 47 12 51
rect 40 47 44 51
rect 58 47 62 51
rect 115 47 119 51
rect 130 47 134 51
rect 158 47 162 51
rect 3 35 7 39
rect 35 33 39 37
rect 55 36 59 40
rect 74 32 78 36
rect 93 33 97 37
rect 112 33 116 37
rect 125 34 129 38
rect 261 59 265 63
rect 283 59 287 63
rect 342 59 346 63
rect 367 59 371 63
rect 398 59 402 63
rect 283 51 287 55
rect 326 52 330 56
rect 348 51 355 55
rect 398 52 402 56
rect 301 47 305 51
rect 319 47 323 51
rect 376 47 380 51
rect 391 47 395 51
rect 419 47 423 51
rect 222 43 226 47
rect 147 33 151 37
rect 155 34 159 38
rect 167 34 171 38
rect 201 28 205 32
rect 241 34 245 38
rect 230 27 234 31
rect 8 17 12 21
rect 33 14 37 18
rect 40 17 44 21
rect 58 17 62 21
rect 80 14 84 18
rect 105 14 109 18
rect 115 17 119 21
rect 131 17 135 21
rect 151 14 155 18
rect 158 17 162 21
rect 296 33 300 37
rect 316 36 320 40
rect 335 32 339 36
rect 354 33 358 37
rect 373 33 377 37
rect 386 34 390 38
rect 408 33 412 37
rect 416 34 420 38
rect 428 34 432 38
rect 242 17 246 21
rect 268 17 272 21
rect 34 7 38 11
rect 65 7 69 11
rect 87 7 91 11
rect 152 7 156 11
rect 294 14 298 18
rect 301 17 305 21
rect 319 17 323 21
rect 341 14 345 18
rect 366 14 370 18
rect 376 17 380 21
rect 392 17 396 21
rect 412 14 416 18
rect 419 17 423 21
rect 212 7 216 11
rect 251 7 255 11
rect 295 7 299 11
rect 326 7 330 11
rect 348 7 352 11
rect 413 7 417 11
rect 7 0 11 4
rect 41 0 45 4
rect 58 0 62 4
rect 114 0 118 4
rect 131 0 135 4
rect 159 0 163 4
rect 242 0 246 4
rect 268 0 272 4
rect 302 0 306 4
rect 319 0 323 4
rect 375 0 379 4
rect 392 0 396 4
rect 420 0 424 4
rect 250 -17 254 -13
rect -30 -25 -26 -21
rect 260 -24 264 -20
<< metal2 >>
rect 10 602 13 612
rect 0 578 3 581
rect 17 572 20 581
rect 33 574 36 587
rect 46 559 49 612
rect 113 602 116 612
rect 142 602 145 612
rect 53 587 57 591
rect 54 572 57 581
rect 9 545 12 557
rect 50 555 51 559
rect 60 545 63 598
rect 66 578 69 583
rect 75 572 78 581
rect 91 574 94 587
rect 112 572 115 581
rect 128 581 131 583
rect 128 578 135 581
rect 128 572 131 578
rect 149 572 152 581
rect 165 574 168 587
rect 111 545 114 555
rect -53 541 -4 545
rect 128 538 131 568
rect 178 559 181 612
rect 245 602 248 612
rect 274 602 277 612
rect 185 587 189 591
rect 186 572 189 581
rect 141 545 144 557
rect 182 555 183 559
rect 192 545 195 598
rect 198 578 201 583
rect 207 572 210 581
rect 223 574 226 587
rect 244 572 247 581
rect 260 581 263 583
rect 260 578 267 581
rect 260 572 263 578
rect 281 572 284 581
rect 297 574 300 587
rect 243 545 246 555
rect 128 535 180 538
rect 8 515 11 528
rect 34 518 37 521
rect 41 515 44 528
rect 58 515 61 528
rect -53 469 -3 473
rect 8 466 11 481
rect 22 473 25 477
rect 40 466 43 481
rect 59 466 62 481
rect 65 480 68 521
rect 81 473 84 514
rect 87 481 90 521
rect 106 473 109 514
rect 115 515 118 528
rect 131 515 134 528
rect 152 518 155 521
rect 159 515 162 528
rect 177 524 180 535
rect 260 532 263 568
rect 310 559 313 612
rect 377 602 380 612
rect 406 602 409 612
rect 317 587 321 591
rect 318 572 321 581
rect 273 545 276 557
rect 314 555 315 559
rect 324 545 327 598
rect 330 578 333 583
rect 339 572 342 581
rect 355 574 358 587
rect 376 572 379 581
rect 392 581 395 583
rect 392 578 399 581
rect 392 572 395 578
rect 413 572 416 581
rect 429 574 432 587
rect 375 545 378 555
rect 392 538 395 560
rect 442 559 445 612
rect 509 602 512 612
rect 449 587 453 591
rect 450 572 453 581
rect 405 545 408 557
rect 446 555 447 559
rect 456 545 459 598
rect 462 578 465 583
rect 471 572 474 581
rect 487 574 490 587
rect 508 572 511 581
rect 524 581 527 583
rect 524 578 528 581
rect 524 572 527 578
rect 507 545 510 555
rect 258 527 263 532
rect 320 534 395 538
rect 177 521 222 524
rect 177 511 180 521
rect 195 508 215 511
rect 212 489 215 508
rect 115 466 118 481
rect 130 466 133 481
rect 137 473 141 476
rect 158 466 161 481
rect -53 455 -3 459
rect 8 447 11 462
rect 22 451 25 455
rect 40 447 43 462
rect 59 447 62 462
rect 8 400 11 413
rect 34 407 37 410
rect 8 383 11 396
rect 41 400 44 413
rect 58 400 61 413
rect 65 407 68 448
rect 81 414 84 455
rect 87 407 90 447
rect 106 414 109 455
rect 115 447 118 462
rect 130 447 133 462
rect 137 452 141 455
rect 158 447 161 462
rect 115 400 118 413
rect 34 386 37 389
rect 41 383 44 396
rect 58 383 61 396
rect -53 337 -3 341
rect 8 334 11 349
rect 22 341 25 345
rect 40 334 43 349
rect 59 334 62 349
rect 65 348 68 389
rect 81 341 84 382
rect 87 349 90 389
rect 106 341 109 382
rect 115 383 118 396
rect 131 400 134 413
rect 152 407 155 410
rect 159 400 162 413
rect 212 413 215 485
rect 223 449 226 521
rect 258 524 261 527
rect 258 521 303 524
rect 258 511 261 521
rect 131 383 134 396
rect 152 386 155 389
rect 159 383 162 396
rect 212 379 215 409
rect 223 393 226 445
rect 230 433 234 499
rect 218 389 222 392
rect 211 376 215 379
rect 212 357 215 376
rect 115 334 118 349
rect 130 334 133 349
rect 137 341 141 344
rect 158 334 161 349
rect -53 323 -3 327
rect 1 323 3 327
rect 8 315 11 330
rect 22 319 25 323
rect 40 315 43 330
rect 59 315 62 330
rect 8 268 11 281
rect 34 275 37 278
rect 8 251 11 264
rect 41 268 44 281
rect 58 268 61 281
rect 65 275 68 316
rect 81 282 84 323
rect 87 275 90 315
rect 106 282 109 323
rect 115 315 118 330
rect 130 315 133 330
rect 137 320 141 323
rect 158 315 161 330
rect 115 268 118 281
rect 34 254 37 257
rect 41 251 44 264
rect 58 251 61 264
rect -53 205 -3 209
rect 8 202 11 217
rect 22 209 25 213
rect 40 202 43 217
rect 59 202 62 217
rect 65 216 68 257
rect 81 209 84 250
rect 87 217 90 257
rect 106 209 109 250
rect 115 251 118 264
rect 131 268 134 281
rect 152 275 155 278
rect 159 268 162 281
rect 212 282 215 353
rect 223 318 226 389
rect 131 251 134 264
rect 152 254 155 257
rect 159 251 162 264
rect 212 225 215 278
rect 223 261 226 314
rect 230 302 234 367
rect 218 257 222 260
rect 261 260 264 511
rect 276 508 296 511
rect 293 489 296 508
rect 293 413 296 485
rect 304 449 307 521
rect 311 433 315 499
rect 320 400 323 534
rect 524 531 527 560
rect 348 528 527 531
rect 282 396 323 400
rect 282 392 285 396
rect 282 389 327 392
rect 282 379 285 389
rect 300 376 320 379
rect 282 374 285 375
rect 317 357 320 376
rect 317 282 320 353
rect 328 318 331 389
rect 335 302 339 367
rect 115 202 118 217
rect 130 202 133 217
rect 137 209 141 212
rect 158 202 161 217
rect -53 191 -3 195
rect 8 183 11 198
rect 22 187 25 191
rect 40 183 43 198
rect 59 183 62 198
rect 8 136 11 149
rect 34 143 37 146
rect 8 119 11 132
rect 41 136 44 149
rect 58 136 61 149
rect 65 143 68 184
rect 81 150 84 191
rect 87 143 90 183
rect 106 150 109 191
rect 115 183 118 198
rect 130 183 133 198
rect 137 188 141 191
rect 158 183 161 198
rect 115 136 118 149
rect 34 122 37 125
rect 41 119 44 132
rect 58 119 61 132
rect -53 73 -3 77
rect 8 70 11 85
rect 22 77 25 81
rect 40 70 43 85
rect 59 70 62 85
rect 65 84 68 125
rect 81 77 84 118
rect 87 85 90 125
rect 106 77 109 118
rect 115 119 118 132
rect 131 136 134 149
rect 152 143 155 146
rect 159 136 162 149
rect 212 147 215 221
rect 223 183 226 257
rect 258 257 303 260
rect 258 247 261 257
rect 276 244 296 247
rect 131 119 134 132
rect 152 122 155 125
rect 159 119 162 132
rect 212 93 215 143
rect 223 129 226 179
rect 230 167 234 235
rect 293 225 296 244
rect 293 147 296 221
rect 304 183 307 257
rect 348 260 351 528
rect 348 257 393 260
rect 348 247 351 257
rect 366 244 386 247
rect 311 167 315 235
rect 383 225 386 244
rect 383 147 386 221
rect 394 183 397 257
rect 401 167 405 235
rect 218 125 222 128
rect 115 70 118 85
rect 130 70 133 85
rect 137 77 141 80
rect 158 70 161 85
rect -53 59 -3 63
rect 8 51 11 66
rect 22 55 25 59
rect 40 51 43 66
rect 59 51 62 66
rect 8 4 11 17
rect 34 11 37 14
rect 41 4 44 17
rect 58 4 61 17
rect 65 11 68 52
rect 81 18 84 59
rect 87 11 90 51
rect 106 18 109 59
rect 115 51 118 66
rect 130 51 133 66
rect 137 56 141 59
rect 158 51 161 66
rect 115 4 118 17
rect 131 4 134 17
rect 152 11 155 14
rect 159 4 162 17
rect 212 11 215 89
rect 223 47 226 125
rect 230 31 234 103
rect 242 4 246 17
rect 251 -13 254 7
rect 261 -20 264 59
rect 283 55 286 59
rect 301 51 304 66
rect 320 51 323 66
rect 268 4 272 17
rect 295 11 298 14
rect 302 4 305 17
rect 319 4 322 17
rect 326 11 329 52
rect 342 18 345 59
rect 348 11 351 51
rect 367 18 370 59
rect 376 51 379 66
rect 391 51 394 66
rect 398 56 402 59
rect 419 51 422 66
rect 376 4 379 17
rect 392 4 395 17
rect 413 11 416 14
rect 420 4 423 17
rect -53 -25 -30 -21
<< m3contact >>
rect 2 498 7 503
rect 39 495 44 500
rect 50 491 55 496
rect 73 500 78 505
rect 97 495 102 500
rect 112 499 117 505
rect 142 495 147 500
rect 171 494 176 499
rect 126 489 131 494
rect 155 489 159 494
rect 197 488 202 493
rect 3 435 8 440
rect 39 428 44 433
rect 50 432 55 437
rect 73 423 78 428
rect 97 428 102 433
rect 126 434 131 439
rect 155 434 159 439
rect 112 423 117 429
rect 142 428 147 433
rect 171 429 176 434
rect 197 429 202 434
rect 2 366 7 371
rect 39 363 44 368
rect 50 359 55 364
rect 73 368 78 373
rect 97 363 102 368
rect 253 494 258 499
rect 112 367 117 373
rect 142 363 147 368
rect 171 362 176 367
rect 126 357 131 362
rect 155 357 159 362
rect 197 356 202 361
rect 3 303 8 308
rect 39 296 44 301
rect 50 300 55 305
rect 73 291 78 296
rect 97 296 102 301
rect 126 302 131 307
rect 155 302 159 307
rect 112 291 117 297
rect 142 296 147 301
rect 171 297 176 302
rect 196 298 201 303
rect 2 234 7 239
rect 39 231 44 236
rect 50 227 55 232
rect 73 236 78 241
rect 97 231 102 236
rect 112 235 117 241
rect 142 231 147 236
rect 171 230 176 235
rect 126 225 131 230
rect 155 225 159 230
rect 197 224 202 229
rect 253 370 258 375
rect 278 488 283 493
rect 277 429 282 434
rect 338 494 343 499
rect 302 356 307 361
rect 302 298 307 303
rect 3 171 8 176
rect 39 164 44 169
rect 50 168 55 173
rect 73 159 78 164
rect 97 164 102 169
rect 126 170 131 175
rect 155 170 159 175
rect 112 159 117 165
rect 142 164 147 169
rect 171 165 176 170
rect 197 163 202 168
rect 2 102 7 107
rect 39 99 44 104
rect 50 95 55 100
rect 73 104 78 109
rect 97 99 102 104
rect 112 103 117 109
rect 142 99 147 104
rect 171 98 176 103
rect 126 93 131 98
rect 155 93 159 98
rect 197 92 202 97
rect 253 230 258 235
rect 278 224 283 229
rect 277 163 282 168
rect 360 367 365 372
rect 335 239 340 244
rect 369 232 374 237
rect 366 159 371 164
rect 425 242 430 247
rect 3 39 8 44
rect 39 32 44 37
rect 50 36 55 41
rect 73 27 78 32
rect 97 32 102 37
rect 126 38 131 43
rect 155 38 159 43
rect 112 27 117 33
rect 142 32 147 37
rect 171 33 176 38
rect 196 27 201 32
rect 253 106 258 111
rect 241 38 246 43
rect 300 32 305 37
rect 311 36 316 41
rect 334 27 339 32
rect 358 32 363 37
rect 387 38 392 43
rect 416 38 420 43
rect 373 27 378 33
rect 403 32 408 37
rect 428 38 433 43
<< metal3 >>
rect 39 505 79 506
rect 1 503 8 504
rect 1 498 2 503
rect 7 498 8 503
rect 39 501 73 505
rect 1 497 8 498
rect 38 500 45 501
rect 38 495 39 500
rect 44 495 45 500
rect 72 500 73 501
rect 78 500 79 505
rect 111 505 147 510
rect 72 499 79 500
rect 96 500 103 501
rect 38 494 45 495
rect 49 496 56 497
rect 49 491 50 496
rect 55 491 56 496
rect 96 495 97 500
rect 102 495 103 500
rect 111 499 112 505
rect 117 504 147 505
rect 117 499 118 504
rect 142 501 147 504
rect 111 498 118 499
rect 141 500 148 501
rect 141 495 142 500
rect 147 495 148 500
rect 170 499 177 500
rect 96 494 103 495
rect 125 494 132 495
rect 141 494 148 495
rect 154 494 160 495
rect 97 491 102 494
rect 49 486 102 491
rect 125 489 126 494
rect 131 489 132 494
rect 154 489 155 494
rect 159 489 160 494
rect 125 488 160 489
rect 126 484 160 488
rect 170 494 171 499
rect 176 494 177 499
rect 252 499 259 500
rect 252 494 253 499
rect 258 494 259 499
rect 337 499 344 500
rect 337 494 338 499
rect 343 494 344 499
rect 170 493 177 494
rect 196 493 203 494
rect 252 493 259 494
rect 277 493 284 494
rect 337 493 344 494
rect 170 488 197 493
rect 202 488 203 493
rect 253 488 278 493
rect 283 488 284 493
rect 170 467 175 488
rect 196 487 203 488
rect 277 487 284 488
rect 334 488 343 493
rect 3 461 175 467
rect 3 441 8 461
rect 2 440 9 441
rect 2 435 3 440
rect 8 435 9 440
rect 2 434 9 435
rect 49 437 102 442
rect 126 440 160 444
rect 38 433 45 434
rect 38 428 39 433
rect 44 428 45 433
rect 49 432 50 437
rect 55 432 56 437
rect 97 434 102 437
rect 125 439 160 440
rect 125 434 126 439
rect 131 434 132 439
rect 154 434 155 439
rect 159 434 160 439
rect 49 431 56 432
rect 96 433 103 434
rect 125 433 132 434
rect 141 433 148 434
rect 154 433 160 434
rect 170 434 177 435
rect 196 434 203 435
rect 276 434 283 435
rect 38 427 45 428
rect 72 428 79 429
rect 72 427 73 428
rect 39 423 73 427
rect 78 423 79 428
rect 96 428 97 433
rect 102 428 103 433
rect 96 427 103 428
rect 111 429 118 430
rect 39 422 79 423
rect 111 423 112 429
rect 117 424 118 429
rect 141 428 142 433
rect 147 428 148 433
rect 170 429 171 434
rect 176 429 197 434
rect 202 429 203 434
rect 170 428 177 429
rect 196 428 203 429
rect 253 429 277 434
rect 282 429 283 434
rect 141 427 148 428
rect 142 424 147 427
rect 117 423 147 424
rect 111 418 147 423
rect 171 401 176 428
rect 2 395 176 401
rect 2 372 7 395
rect 39 373 79 374
rect 1 371 8 372
rect 1 366 2 371
rect 7 366 8 371
rect 39 369 73 373
rect 1 365 8 366
rect 38 368 45 369
rect 38 363 39 368
rect 44 363 45 368
rect 72 368 73 369
rect 78 368 79 373
rect 111 373 147 378
rect 253 376 258 429
rect 276 428 283 429
rect 334 400 339 488
rect 296 395 339 400
rect 72 367 79 368
rect 96 368 103 369
rect 38 362 45 363
rect 49 364 56 365
rect 49 359 50 364
rect 55 359 56 364
rect 96 363 97 368
rect 102 363 103 368
rect 111 367 112 373
rect 117 372 147 373
rect 117 367 118 372
rect 142 369 147 372
rect 252 375 259 376
rect 252 370 253 375
rect 258 370 259 375
rect 252 369 259 370
rect 111 366 118 367
rect 141 368 148 369
rect 141 363 142 368
rect 147 363 148 368
rect 170 367 177 368
rect 96 362 103 363
rect 125 362 132 363
rect 141 362 148 363
rect 154 362 160 363
rect 97 359 102 362
rect 49 354 102 359
rect 125 357 126 362
rect 131 357 132 362
rect 154 357 155 362
rect 159 357 160 362
rect 125 356 160 357
rect 126 352 160 356
rect 170 362 171 367
rect 176 362 177 367
rect 296 362 301 395
rect 359 372 366 373
rect 359 367 360 372
rect 365 367 366 372
rect 359 366 366 367
rect 170 361 177 362
rect 196 361 203 362
rect 170 356 197 361
rect 202 356 203 361
rect 296 361 308 362
rect 296 356 302 361
rect 307 356 308 361
rect 170 335 175 356
rect 196 355 203 356
rect 301 355 308 356
rect 3 329 175 335
rect 3 309 8 329
rect 2 308 9 309
rect 2 303 3 308
rect 8 303 9 308
rect 2 302 9 303
rect 49 305 102 310
rect 126 308 160 312
rect 38 301 45 302
rect 38 296 39 301
rect 44 296 45 301
rect 49 300 50 305
rect 55 300 56 305
rect 97 302 102 305
rect 125 307 160 308
rect 125 302 126 307
rect 131 302 132 307
rect 154 302 155 307
rect 159 302 160 307
rect 195 303 202 304
rect 301 303 308 304
rect 49 299 56 300
rect 96 301 103 302
rect 125 301 132 302
rect 141 301 148 302
rect 154 301 160 302
rect 170 302 196 303
rect 38 295 45 296
rect 72 296 79 297
rect 72 295 73 296
rect 39 291 73 295
rect 78 291 79 296
rect 96 296 97 301
rect 102 296 103 301
rect 96 295 103 296
rect 111 297 118 298
rect 39 290 79 291
rect 111 291 112 297
rect 117 292 118 297
rect 141 296 142 301
rect 147 296 148 301
rect 141 295 148 296
rect 170 297 171 302
rect 176 298 196 302
rect 201 298 202 303
rect 176 297 177 298
rect 195 297 202 298
rect 297 298 302 303
rect 307 298 308 303
rect 297 297 308 298
rect 170 296 177 297
rect 142 292 147 295
rect 117 291 147 292
rect 111 286 147 291
rect 170 269 175 296
rect 2 263 175 269
rect 297 269 302 297
rect 297 264 340 269
rect 2 240 7 263
rect 39 241 79 242
rect 1 239 8 240
rect 1 234 2 239
rect 7 234 8 239
rect 39 237 73 241
rect 1 233 8 234
rect 38 236 45 237
rect 38 231 39 236
rect 44 231 45 236
rect 72 236 73 237
rect 78 236 79 241
rect 111 241 147 246
rect 335 245 340 264
rect 72 235 79 236
rect 96 236 103 237
rect 38 230 45 231
rect 49 232 56 233
rect 49 227 50 232
rect 55 227 56 232
rect 96 231 97 236
rect 102 231 103 236
rect 111 235 112 241
rect 117 240 147 241
rect 117 235 118 240
rect 142 237 147 240
rect 334 244 341 245
rect 334 239 335 244
rect 340 239 341 244
rect 334 238 341 239
rect 360 237 365 366
rect 424 247 431 248
rect 424 242 425 247
rect 430 242 532 247
rect 424 241 431 242
rect 368 237 375 238
rect 111 234 118 235
rect 141 236 148 237
rect 141 231 142 236
rect 147 231 148 236
rect 170 235 177 236
rect 96 230 103 231
rect 125 230 132 231
rect 141 230 148 231
rect 154 230 160 231
rect 97 227 102 230
rect 49 222 102 227
rect 125 225 126 230
rect 131 225 132 230
rect 154 225 155 230
rect 159 225 160 230
rect 125 224 160 225
rect 126 220 160 224
rect 170 230 171 235
rect 176 230 177 235
rect 252 235 259 236
rect 252 230 253 235
rect 258 230 259 235
rect 348 232 369 237
rect 374 232 375 237
rect 348 231 360 232
rect 368 231 375 232
rect 170 229 177 230
rect 196 229 203 230
rect 252 229 259 230
rect 277 229 284 230
rect 170 224 197 229
rect 202 224 203 229
rect 253 224 278 229
rect 283 224 284 229
rect 170 203 175 224
rect 196 223 203 224
rect 277 223 284 224
rect 348 223 353 231
rect 3 197 175 203
rect 315 202 353 223
rect 3 177 8 197
rect 2 176 9 177
rect 2 171 3 176
rect 8 171 9 176
rect 2 170 9 171
rect 49 173 102 178
rect 126 176 160 180
rect 38 169 45 170
rect 38 164 39 169
rect 44 164 45 169
rect 49 168 50 173
rect 55 168 56 173
rect 97 170 102 173
rect 125 175 160 176
rect 125 170 126 175
rect 131 170 132 175
rect 154 170 155 175
rect 159 170 160 175
rect 49 167 56 168
rect 96 169 103 170
rect 125 169 132 170
rect 141 169 148 170
rect 154 169 160 170
rect 170 170 177 171
rect 38 163 45 164
rect 72 164 79 165
rect 72 163 73 164
rect 39 159 73 163
rect 78 159 79 164
rect 96 164 97 169
rect 102 164 103 169
rect 96 163 103 164
rect 111 165 118 166
rect 39 158 79 159
rect 111 159 112 165
rect 117 160 118 165
rect 141 164 142 169
rect 147 164 148 169
rect 170 165 171 170
rect 176 168 177 170
rect 196 168 203 169
rect 276 168 283 169
rect 176 165 197 168
rect 170 164 197 165
rect 141 163 148 164
rect 171 163 197 164
rect 202 163 203 168
rect 142 160 147 163
rect 117 159 147 160
rect 111 154 147 159
rect 171 137 176 163
rect 196 162 203 163
rect 253 163 277 168
rect 282 163 283 168
rect 2 131 176 137
rect 2 108 7 131
rect 39 109 79 110
rect 1 107 8 108
rect 1 102 2 107
rect 7 102 8 107
rect 39 105 73 109
rect 1 101 8 102
rect 38 104 45 105
rect 38 99 39 104
rect 44 99 45 104
rect 72 104 73 105
rect 78 104 79 109
rect 111 109 147 114
rect 253 112 258 163
rect 276 162 283 163
rect 72 103 79 104
rect 96 104 103 105
rect 38 98 45 99
rect 49 100 56 101
rect 49 95 50 100
rect 55 95 56 100
rect 96 99 97 104
rect 102 99 103 104
rect 111 103 112 109
rect 117 108 147 109
rect 117 103 118 108
rect 142 105 147 108
rect 252 111 259 112
rect 252 106 253 111
rect 258 106 259 111
rect 252 105 259 106
rect 111 102 118 103
rect 141 104 148 105
rect 141 99 142 104
rect 147 99 148 104
rect 170 103 177 104
rect 96 98 103 99
rect 125 98 132 99
rect 141 98 148 99
rect 154 98 160 99
rect 97 95 102 98
rect 49 90 102 95
rect 125 93 126 98
rect 131 93 132 98
rect 154 93 155 98
rect 159 93 160 98
rect 125 92 160 93
rect 126 88 160 92
rect 170 98 171 103
rect 176 98 177 103
rect 170 97 177 98
rect 196 97 203 98
rect 170 92 197 97
rect 202 92 203 97
rect 315 93 320 202
rect 365 164 372 165
rect 365 159 366 164
rect 371 159 372 164
rect 365 158 372 159
rect 272 92 320 93
rect 170 71 175 92
rect 196 91 203 92
rect 3 65 175 71
rect 241 87 320 92
rect 366 96 371 158
rect 366 90 433 96
rect 3 45 8 65
rect 2 44 9 45
rect 2 39 3 44
rect 8 39 9 44
rect 2 38 9 39
rect 49 41 102 46
rect 126 44 160 48
rect 241 44 246 87
rect 38 37 45 38
rect 38 32 39 37
rect 44 32 45 37
rect 49 36 50 41
rect 55 36 56 41
rect 97 38 102 41
rect 125 43 160 44
rect 125 38 126 43
rect 131 38 132 43
rect 154 38 155 43
rect 159 38 160 43
rect 240 43 247 44
rect 49 35 56 36
rect 96 37 103 38
rect 125 37 132 38
rect 141 37 148 38
rect 154 37 160 38
rect 170 38 177 39
rect 38 31 45 32
rect 72 32 79 33
rect 72 31 73 32
rect 39 27 73 31
rect 78 27 79 32
rect 96 32 97 37
rect 102 32 103 37
rect 96 31 103 32
rect 111 33 118 34
rect 39 26 79 27
rect 111 27 112 33
rect 117 28 118 33
rect 141 32 142 37
rect 147 32 148 37
rect 170 33 171 38
rect 176 33 177 38
rect 240 38 241 43
rect 246 38 247 43
rect 310 41 363 46
rect 387 44 421 48
rect 428 44 433 90
rect 240 37 247 38
rect 299 37 306 38
rect 170 32 177 33
rect 195 32 202 33
rect 141 31 148 32
rect 142 28 147 31
rect 117 27 147 28
rect 172 27 196 32
rect 201 27 202 32
rect 299 32 300 37
rect 305 32 306 37
rect 310 36 311 41
rect 316 36 317 41
rect 358 38 363 41
rect 386 43 421 44
rect 386 38 387 43
rect 392 38 393 43
rect 415 38 416 43
rect 420 38 421 43
rect 310 35 317 36
rect 357 37 364 38
rect 386 37 393 38
rect 402 37 409 38
rect 415 37 421 38
rect 427 43 434 44
rect 427 38 428 43
rect 433 38 434 43
rect 427 37 434 38
rect 299 31 306 32
rect 333 32 340 33
rect 333 31 334 32
rect 111 22 147 27
rect 195 26 202 27
rect 300 27 334 31
rect 339 27 340 32
rect 357 32 358 37
rect 363 32 364 37
rect 357 31 364 32
rect 372 33 379 34
rect 300 26 340 27
rect 372 27 373 33
rect 378 28 379 33
rect 402 32 403 37
rect 408 32 409 37
rect 402 31 409 32
rect 403 28 408 31
rect 378 27 408 28
rect 372 22 408 27
<< labels >>
rlabel metal1 1 521 5 525 3 clk
rlabel metal1 1 528 5 532 3 Vdd!
rlabel metal1 1 469 5 473 3 ~clk
rlabel metal1 1 403 5 407 3 clk
rlabel metal1 1 455 5 459 3 ~clk
rlabel metal1 1 462 5 466 3 GND!
rlabel metal1 1 389 5 393 3 clk
rlabel metal1 1 396 5 400 3 Vdd!
rlabel metal1 1 337 5 341 3 ~clk
rlabel metal1 1 271 5 275 3 clk
rlabel metal1 1 323 5 327 3 ~clk
rlabel metal1 1 330 5 334 3 GND!
rlabel metal1 1 66 5 70 3 GND!
rlabel metal1 1 59 5 63 3 ~clk
rlabel metal1 1 0 5 4 3 Vdd!
rlabel metal1 1 7 5 11 3 clk
rlabel metal1 1 73 5 77 3 ~clk
rlabel metal1 1 132 5 136 3 Vdd!
rlabel metal1 1 125 5 129 3 clk
rlabel metal1 1 198 5 202 3 GND!
rlabel metal1 1 191 5 195 3 ~clk
rlabel metal1 1 139 5 143 3 clk
rlabel metal1 1 205 5 209 3 ~clk
rlabel metal1 1 264 5 268 3 Vdd!
rlabel metal1 1 257 5 261 3 clk
rlabel polysilicon 265 39 267 42 5 reset
rlabel polysilicon 247 30 249 33 5 D
rlabel metal1 203 0 207 4 1 Vdd!
rlabel metal1 204 66 207 70 1 GND!
rlabel metal1 374 132 378 136 1 Vdd!
rlabel metal1 284 132 288 136 1 Vdd!
rlabel metal1 203 132 207 136 1 Vdd!
rlabel metal1 375 198 378 202 1 GND!
rlabel metal1 285 198 288 202 1 GND!
rlabel metal1 204 198 207 202 1 GND!
rlabel metal1 425 235 428 238 7 out
rlabel metal1 374 264 378 268 1 Vdd!
rlabel metal1 203 264 207 268 1 Vdd!
rlabel metal1 284 264 288 268 1 Vdd!
rlabel metal1 204 330 207 334 1 GND!
rlabel metal1 309 330 312 334 1 GND!
rlabel metal1 203 396 207 400 1 Vdd!
rlabel metal1 284 396 288 400 1 Vdd!
rlabel metal1 353 367 356 370 7 Y
rlabel metal1 203 528 207 532 1 Vdd!
rlabel metal1 284 528 288 532 1 Vdd!
rlabel metal1 204 462 207 466 1 GND!
rlabel metal1 285 462 288 466 1 GND!
rlabel metal2 348 523 351 528 1 select_out
rlabel metal1 3 605 6 609 1 Vdd!
rlabel metal1 4 548 7 552 1 GND!
rlabel metal1 5 541 8 545 2 ~clk
rlabel metal1 3 612 6 616 4 clk
rlabel metal1 136 548 139 552 1 GND!
rlabel metal1 137 541 140 545 2 ~clk
rlabel metal1 135 612 138 616 4 clk
rlabel metal1 267 605 270 609 1 Vdd!
rlabel metal1 268 548 271 552 1 GND!
rlabel metal1 269 541 272 545 2 ~clk
rlabel metal1 267 612 270 616 4 clk
rlabel metal1 399 612 402 616 4 clk
rlabel metal1 401 541 404 545 2 ~clk
rlabel metal1 400 548 403 552 1 GND!
rlabel metal1 399 605 402 609 1 Vdd!
rlabel metal2 0 578 3 581 3 ctrl_reg
rlabel metal2 177 533 180 538 1 select0
rlabel metal2 260 532 263 539 1 select1
rlabel metal2 320 532 323 538 1 select2
rlabel m3contact 2 498 7 503 3 data_reg
rlabel metal1 264 0 268 4 1 Vdd!
rlabel metal1 253 66 257 70 1 GND!
rlabel metal1 254 59 258 63 1 ~clk
rlabel metal1 257 7 260 11 1 clk
rlabel metal1 135 605 138 609 1 Vdd!
<< end >>
