magic
tech scmos
timestamp 1608311150
<< ntransistor >>
rect 662 927 664 931
rect 667 927 669 931
rect 683 927 685 931
rect 699 927 701 931
rect 704 927 706 931
rect 725 927 727 931
rect 741 927 743 931
rect 757 927 759 931
rect 762 927 764 931
rect 778 927 780 931
rect 794 927 796 931
rect 799 927 801 931
rect 815 927 817 931
rect 831 927 833 931
rect 836 927 838 931
rect 857 927 859 931
rect 873 927 875 931
rect 889 927 891 931
rect 894 927 896 931
rect 910 927 912 931
rect 926 927 928 931
rect 931 927 933 931
rect 947 927 949 931
rect 963 927 965 931
rect 968 927 970 931
rect 989 927 991 931
rect 1005 927 1007 931
rect 1021 927 1023 931
rect 1026 927 1028 931
rect 1042 927 1044 931
rect 1058 927 1060 931
rect 1063 927 1065 931
rect 1079 927 1081 931
rect 1095 927 1097 931
rect 1100 927 1102 931
rect 1121 927 1123 931
rect 1137 927 1139 931
rect 1153 927 1155 931
rect 1158 927 1160 931
rect 1174 927 1176 931
rect 322 894 324 898
rect 327 894 329 898
rect 343 894 345 898
rect 359 894 361 898
rect 364 894 366 898
rect 385 894 387 898
rect 401 894 403 898
rect 417 894 419 898
rect 422 894 424 898
rect 438 894 440 898
rect 446 857 448 861
rect 841 861 843 865
rect 867 857 869 861
rect 872 857 874 861
rect 922 861 924 865
rect 948 857 950 861
rect 953 857 955 861
rect 895 853 897 857
rect 329 848 331 852
rect 667 848 669 852
rect 683 848 685 852
rect 699 848 701 852
rect 722 848 724 852
rect 727 848 729 852
rect 753 848 755 852
rect 774 848 776 852
rect 794 848 796 852
rect 799 848 801 852
rect 817 848 819 852
rect 976 853 978 857
rect 667 802 669 806
rect 683 802 685 806
rect 699 802 701 806
rect 722 802 724 806
rect 727 802 729 806
rect 753 802 755 806
rect 774 802 776 806
rect 794 802 796 806
rect 799 802 801 806
rect 817 802 819 806
rect 313 792 315 796
rect 329 792 331 796
rect 334 792 336 796
rect 350 792 352 796
rect 366 792 368 796
rect 387 792 389 796
rect 392 792 394 796
rect 408 792 410 796
rect 424 792 426 796
rect 429 792 431 796
rect 867 801 869 805
rect 872 801 874 805
rect 948 801 950 805
rect 953 801 955 805
rect 867 725 869 729
rect 872 725 874 729
rect 946 729 948 733
rect 972 725 974 729
rect 977 725 979 729
rect 895 721 897 725
rect 667 716 669 720
rect 683 716 685 720
rect 699 716 701 720
rect 722 716 724 720
rect 727 716 729 720
rect 753 716 755 720
rect 774 716 776 720
rect 794 716 796 720
rect 799 716 801 720
rect 817 716 819 720
rect 1000 721 1002 725
rect 667 670 669 674
rect 683 670 685 674
rect 699 670 701 674
rect 722 670 724 674
rect 727 670 729 674
rect 753 670 755 674
rect 774 670 776 674
rect 794 670 796 674
rect 799 670 801 674
rect 817 670 819 674
rect 867 670 869 674
rect 872 670 874 674
rect 972 670 974 674
rect 977 670 979 674
rect 867 593 869 597
rect 872 593 874 597
rect 922 597 924 601
rect 948 593 950 597
rect 953 593 955 597
rect 1012 597 1014 601
rect 1038 593 1040 597
rect 1043 593 1045 597
rect 895 589 897 593
rect 667 584 669 588
rect 683 584 685 588
rect 699 584 701 588
rect 722 584 724 588
rect 727 584 729 588
rect 753 584 755 588
rect 774 584 776 588
rect 794 584 796 588
rect 799 584 801 588
rect 817 584 819 588
rect 976 589 978 593
rect 1066 589 1068 593
rect 667 538 669 542
rect 683 538 685 542
rect 699 538 701 542
rect 722 538 724 542
rect 727 538 729 542
rect 753 538 755 542
rect 774 538 776 542
rect 794 538 796 542
rect 799 538 801 542
rect 817 538 819 542
rect 867 535 869 539
rect 872 535 874 539
rect 948 535 950 539
rect 953 535 955 539
rect 1038 535 1040 539
rect 1043 535 1045 539
rect 867 461 869 465
rect 872 461 874 465
rect 895 457 897 461
rect 667 452 669 456
rect 683 452 685 456
rect 699 452 701 456
rect 722 452 724 456
rect 727 452 729 456
rect 753 452 755 456
rect 774 452 776 456
rect 794 452 796 456
rect 799 452 801 456
rect 817 452 819 456
rect 667 406 669 410
rect 683 406 685 410
rect 699 406 701 410
rect 722 406 724 410
rect 727 406 729 410
rect 753 406 755 410
rect 774 406 776 410
rect 794 406 796 410
rect 799 406 801 410
rect 817 406 819 410
rect 901 406 903 410
rect 919 406 921 410
rect 944 406 946 410
rect 960 406 962 410
rect 983 406 985 410
rect 988 406 990 410
rect 1014 406 1016 410
rect 1035 406 1037 410
rect 1055 406 1057 410
rect 1060 406 1062 410
rect 1078 406 1080 410
rect 190 392 192 396
rect 195 392 197 396
rect 211 392 213 396
rect 227 392 229 396
rect 232 392 234 396
rect 253 392 255 396
rect 269 392 271 396
rect 285 392 287 396
rect 290 392 292 396
rect 306 392 308 396
rect 322 392 324 396
rect 327 392 329 396
rect 343 392 345 396
rect 359 392 361 396
rect 364 392 366 396
rect 385 392 387 396
rect 401 392 403 396
rect 417 392 419 396
rect 422 392 424 396
rect 438 392 440 396
rect 454 392 456 396
rect 459 392 461 396
rect 475 392 477 396
rect 491 392 493 396
rect 496 392 498 396
rect 517 392 519 396
rect 533 392 535 396
rect 549 392 551 396
rect 554 392 556 396
rect 570 392 572 396
rect 867 399 869 403
rect 872 399 874 403
rect 305 348 307 352
rect 329 348 331 352
rect 1090 350 1094 352
rect 325 337 327 341
rect 316 323 320 325
rect 305 314 307 318
rect 329 314 331 318
rect 961 282 963 286
rect 966 282 968 286
rect 982 282 984 286
rect 998 282 1000 286
rect 1003 282 1005 286
rect 1024 282 1026 286
rect 1040 282 1042 286
rect 1056 282 1058 286
rect 1061 282 1063 286
rect 1077 282 1079 286
rect 190 252 192 256
rect 195 252 197 256
rect 211 252 213 256
rect 227 252 229 256
rect 232 252 234 256
rect 253 252 255 256
rect 269 252 271 256
rect 285 252 287 256
rect 290 252 292 256
rect 306 252 308 256
rect 322 252 324 256
rect 327 252 329 256
rect 343 252 345 256
rect 359 252 361 256
rect 364 252 366 256
rect 385 252 387 256
rect 401 252 403 256
rect 417 252 419 256
rect 422 252 424 256
rect 438 252 440 256
rect 454 252 456 256
rect 459 252 461 256
rect 475 252 477 256
rect 491 252 493 256
rect 496 252 498 256
rect 517 252 519 256
rect 533 252 535 256
rect 549 252 551 256
rect 554 252 556 256
rect 570 252 572 256
rect 1102 206 1106 208
rect 961 196 963 200
rect 966 196 968 200
rect 982 196 984 200
rect 998 196 1000 200
rect 1003 196 1005 200
rect 1024 196 1026 200
rect 1040 196 1042 200
rect 1056 196 1058 200
rect 1061 196 1063 200
rect 1077 196 1079 200
rect 190 166 192 170
rect 195 166 197 170
rect 211 166 213 170
rect 227 166 229 170
rect 232 166 234 170
rect 253 166 255 170
rect 269 166 271 170
rect 285 166 287 170
rect 290 166 292 170
rect 306 166 308 170
rect 322 166 324 170
rect 327 166 329 170
rect 343 166 345 170
rect 359 166 361 170
rect 364 166 366 170
rect 385 166 387 170
rect 401 166 403 170
rect 417 166 419 170
rect 422 166 424 170
rect 438 166 440 170
rect 454 166 456 170
rect 459 166 461 170
rect 475 166 477 170
rect 491 166 493 170
rect 496 166 498 170
rect 517 166 519 170
rect 533 166 535 170
rect 549 166 551 170
rect 554 166 556 170
rect 570 166 572 170
rect 422 122 424 126
rect 446 122 448 126
rect 442 111 444 115
rect 433 97 437 99
rect 422 88 424 92
rect 446 88 448 92
rect 190 26 192 30
rect 195 26 197 30
rect 211 26 213 30
rect 227 26 229 30
rect 232 26 234 30
rect 253 26 255 30
rect 269 26 271 30
rect 285 26 287 30
rect 290 26 292 30
rect 306 26 308 30
rect 322 26 324 30
rect 327 26 329 30
rect 343 26 345 30
rect 359 26 361 30
rect 364 26 366 30
rect 385 26 387 30
rect 401 26 403 30
rect 417 26 419 30
rect 422 26 424 30
rect 438 26 440 30
rect 454 26 456 30
rect 459 26 461 30
rect 475 26 477 30
rect 491 26 493 30
rect 496 26 498 30
rect 517 26 519 30
rect 533 26 535 30
rect 549 26 551 30
rect 554 26 556 30
rect 570 26 572 30
<< ptransistor >>
rect 662 950 664 958
rect 667 950 669 958
rect 683 950 685 958
rect 699 950 701 958
rect 704 950 706 958
rect 725 950 727 958
rect 741 950 743 958
rect 757 950 759 958
rect 762 950 764 958
rect 778 950 780 958
rect 794 950 796 958
rect 799 950 801 958
rect 815 950 817 958
rect 831 950 833 958
rect 836 950 838 958
rect 857 950 859 958
rect 873 950 875 958
rect 889 950 891 958
rect 894 950 896 958
rect 910 950 912 958
rect 926 950 928 958
rect 931 950 933 958
rect 947 950 949 958
rect 963 950 965 958
rect 968 950 970 958
rect 989 950 991 958
rect 1005 950 1007 958
rect 1021 950 1023 958
rect 1026 950 1028 958
rect 1042 950 1044 958
rect 1058 950 1060 958
rect 1063 950 1065 958
rect 1079 950 1081 958
rect 1095 950 1097 958
rect 1100 950 1102 958
rect 1121 950 1123 958
rect 1137 950 1139 958
rect 1153 950 1155 958
rect 1158 950 1160 958
rect 1174 950 1176 958
rect 322 917 324 925
rect 327 917 329 925
rect 343 917 345 925
rect 359 917 361 925
rect 364 917 366 925
rect 385 917 387 925
rect 401 917 403 925
rect 417 917 419 925
rect 422 917 424 925
rect 438 917 440 925
rect 841 879 843 887
rect 667 866 669 874
rect 683 866 685 874
rect 699 866 701 874
rect 722 866 724 874
rect 727 866 729 874
rect 753 866 755 874
rect 774 866 776 874
rect 794 866 796 874
rect 799 866 801 874
rect 817 866 819 874
rect 867 873 869 881
rect 872 873 874 881
rect 895 879 897 887
rect 922 879 924 887
rect 948 873 950 881
rect 953 873 955 881
rect 976 879 978 887
rect 313 815 315 823
rect 329 815 331 823
rect 334 815 336 823
rect 350 815 352 823
rect 366 815 368 823
rect 387 815 389 823
rect 392 815 394 823
rect 408 815 410 823
rect 424 815 426 823
rect 429 815 431 823
rect 667 780 669 788
rect 683 780 685 788
rect 699 780 701 788
rect 722 780 724 788
rect 727 780 729 788
rect 753 780 755 788
rect 774 780 776 788
rect 794 780 796 788
rect 799 780 801 788
rect 817 780 819 788
rect 867 781 869 789
rect 872 781 874 789
rect 948 781 950 789
rect 953 781 955 789
rect 667 734 669 742
rect 683 734 685 742
rect 699 734 701 742
rect 722 734 724 742
rect 727 734 729 742
rect 753 734 755 742
rect 774 734 776 742
rect 794 734 796 742
rect 799 734 801 742
rect 817 734 819 742
rect 867 741 869 749
rect 872 741 874 749
rect 895 747 897 755
rect 946 747 948 755
rect 972 741 974 749
rect 977 741 979 749
rect 1000 747 1002 755
rect 667 648 669 656
rect 683 648 685 656
rect 699 648 701 656
rect 722 648 724 656
rect 727 648 729 656
rect 753 648 755 656
rect 774 648 776 656
rect 794 648 796 656
rect 799 648 801 656
rect 817 648 819 656
rect 867 650 869 658
rect 872 650 874 658
rect 972 650 974 658
rect 977 650 979 658
rect 667 602 669 610
rect 683 602 685 610
rect 699 602 701 610
rect 722 602 724 610
rect 727 602 729 610
rect 753 602 755 610
rect 774 602 776 610
rect 794 602 796 610
rect 799 602 801 610
rect 817 602 819 610
rect 867 609 869 617
rect 872 609 874 617
rect 895 615 897 623
rect 922 615 924 623
rect 948 609 950 617
rect 953 609 955 617
rect 976 615 978 623
rect 1012 615 1014 623
rect 1038 609 1040 617
rect 1043 609 1045 617
rect 1066 615 1068 623
rect 667 516 669 524
rect 683 516 685 524
rect 699 516 701 524
rect 722 516 724 524
rect 727 516 729 524
rect 753 516 755 524
rect 774 516 776 524
rect 794 516 796 524
rect 799 516 801 524
rect 817 516 819 524
rect 867 515 869 523
rect 872 515 874 523
rect 948 515 950 523
rect 953 515 955 523
rect 1038 515 1040 523
rect 1043 515 1045 523
rect 667 470 669 478
rect 683 470 685 478
rect 699 470 701 478
rect 722 470 724 478
rect 727 470 729 478
rect 753 470 755 478
rect 774 470 776 478
rect 794 470 796 478
rect 799 470 801 478
rect 817 470 819 478
rect 867 477 869 485
rect 872 477 874 485
rect 895 483 897 491
rect 190 415 192 423
rect 195 415 197 423
rect 211 415 213 423
rect 227 415 229 423
rect 232 415 234 423
rect 253 415 255 423
rect 269 415 271 423
rect 285 415 287 423
rect 290 415 292 423
rect 306 415 308 423
rect 322 415 324 423
rect 327 415 329 423
rect 343 415 345 423
rect 359 415 361 423
rect 364 415 366 423
rect 385 415 387 423
rect 401 415 403 423
rect 417 415 419 423
rect 422 415 424 423
rect 438 415 440 423
rect 454 415 456 423
rect 459 415 461 423
rect 475 415 477 423
rect 491 415 493 423
rect 496 415 498 423
rect 517 415 519 423
rect 533 415 535 423
rect 549 415 551 423
rect 554 415 556 423
rect 570 415 572 423
rect 667 384 669 392
rect 683 384 685 392
rect 699 384 701 392
rect 722 384 724 392
rect 727 384 729 392
rect 753 384 755 392
rect 774 384 776 392
rect 794 384 796 392
rect 799 384 801 392
rect 817 384 819 392
rect 867 379 869 387
rect 872 379 874 387
rect 901 384 903 392
rect 919 384 921 392
rect 944 384 946 392
rect 960 384 962 392
rect 983 384 985 392
rect 988 384 990 392
rect 1014 384 1016 392
rect 1035 384 1037 392
rect 1055 384 1057 392
rect 1060 384 1062 392
rect 1078 384 1080 392
rect 961 305 963 313
rect 966 305 968 313
rect 982 305 984 313
rect 998 305 1000 313
rect 1003 305 1005 313
rect 1024 305 1026 313
rect 1040 305 1042 313
rect 1056 305 1058 313
rect 1061 305 1063 313
rect 1077 305 1079 313
rect 190 275 192 283
rect 195 275 197 283
rect 211 275 213 283
rect 227 275 229 283
rect 232 275 234 283
rect 253 275 255 283
rect 269 275 271 283
rect 285 275 287 283
rect 290 275 292 283
rect 306 275 308 283
rect 322 275 324 283
rect 327 275 329 283
rect 343 275 345 283
rect 359 275 361 283
rect 364 275 366 283
rect 385 275 387 283
rect 401 275 403 283
rect 417 275 419 283
rect 422 275 424 283
rect 438 275 440 283
rect 454 275 456 283
rect 459 275 461 283
rect 475 275 477 283
rect 491 275 493 283
rect 496 275 498 283
rect 517 275 519 283
rect 533 275 535 283
rect 549 275 551 283
rect 554 275 556 283
rect 570 275 572 283
rect 961 219 963 227
rect 966 219 968 227
rect 982 219 984 227
rect 998 219 1000 227
rect 1003 219 1005 227
rect 1024 219 1026 227
rect 1040 219 1042 227
rect 1056 219 1058 227
rect 1061 219 1063 227
rect 1077 219 1079 227
rect 190 189 192 197
rect 195 189 197 197
rect 211 189 213 197
rect 227 189 229 197
rect 232 189 234 197
rect 253 189 255 197
rect 269 189 271 197
rect 285 189 287 197
rect 290 189 292 197
rect 306 189 308 197
rect 322 189 324 197
rect 327 189 329 197
rect 343 189 345 197
rect 359 189 361 197
rect 364 189 366 197
rect 385 189 387 197
rect 401 189 403 197
rect 417 189 419 197
rect 422 189 424 197
rect 438 189 440 197
rect 454 189 456 197
rect 459 189 461 197
rect 475 189 477 197
rect 491 189 493 197
rect 496 189 498 197
rect 517 189 519 197
rect 533 189 535 197
rect 549 189 551 197
rect 554 189 556 197
rect 570 189 572 197
rect 190 49 192 57
rect 195 49 197 57
rect 211 49 213 57
rect 227 49 229 57
rect 232 49 234 57
rect 253 49 255 57
rect 269 49 271 57
rect 285 49 287 57
rect 290 49 292 57
rect 306 49 308 57
rect 322 49 324 57
rect 327 49 329 57
rect 343 49 345 57
rect 359 49 361 57
rect 364 49 366 57
rect 385 49 387 57
rect 401 49 403 57
rect 417 49 419 57
rect 422 49 424 57
rect 438 49 440 57
rect 454 49 456 57
rect 459 49 461 57
rect 475 49 477 57
rect 491 49 493 57
rect 496 49 498 57
rect 517 49 519 57
rect 533 49 535 57
rect 549 49 551 57
rect 554 49 556 57
rect 570 49 572 57
<< ndiffusion >>
rect 661 927 662 931
rect 664 927 667 931
rect 669 927 670 931
rect 682 927 683 931
rect 685 927 686 931
rect 698 927 699 931
rect 701 927 704 931
rect 706 927 707 931
rect 724 927 725 931
rect 727 927 728 931
rect 740 927 741 931
rect 743 927 744 931
rect 756 927 757 931
rect 759 927 762 931
rect 764 927 765 931
rect 777 927 778 931
rect 780 927 781 931
rect 793 927 794 931
rect 796 927 799 931
rect 801 927 802 931
rect 814 927 815 931
rect 817 927 818 931
rect 830 927 831 931
rect 833 927 836 931
rect 838 927 839 931
rect 856 927 857 931
rect 859 927 860 931
rect 872 927 873 931
rect 875 927 876 931
rect 888 927 889 931
rect 891 927 894 931
rect 896 927 897 931
rect 909 927 910 931
rect 912 927 913 931
rect 925 927 926 931
rect 928 927 931 931
rect 933 927 934 931
rect 946 927 947 931
rect 949 927 950 931
rect 962 927 963 931
rect 965 927 968 931
rect 970 927 971 931
rect 988 927 989 931
rect 991 927 992 931
rect 1004 927 1005 931
rect 1007 927 1008 931
rect 1020 927 1021 931
rect 1023 927 1026 931
rect 1028 927 1029 931
rect 1041 927 1042 931
rect 1044 927 1045 931
rect 1057 927 1058 931
rect 1060 927 1063 931
rect 1065 927 1066 931
rect 1078 927 1079 931
rect 1081 927 1082 931
rect 1094 927 1095 931
rect 1097 927 1100 931
rect 1102 927 1103 931
rect 1120 927 1121 931
rect 1123 927 1124 931
rect 1136 927 1137 931
rect 1139 927 1140 931
rect 1152 927 1153 931
rect 1155 927 1158 931
rect 1160 927 1161 931
rect 1173 927 1174 931
rect 1176 927 1177 931
rect 321 894 322 898
rect 324 894 327 898
rect 329 894 330 898
rect 342 894 343 898
rect 345 894 346 898
rect 358 894 359 898
rect 361 894 364 898
rect 366 894 367 898
rect 384 894 385 898
rect 387 894 388 898
rect 400 894 401 898
rect 403 894 404 898
rect 416 894 417 898
rect 419 894 422 898
rect 424 894 425 898
rect 437 894 438 898
rect 440 894 441 898
rect 445 857 446 861
rect 448 857 449 861
rect 840 861 841 865
rect 843 861 844 865
rect 864 857 867 861
rect 869 857 872 861
rect 874 857 875 861
rect 921 861 922 865
rect 924 861 925 865
rect 945 857 948 861
rect 950 857 953 861
rect 955 857 956 861
rect 894 853 895 857
rect 897 853 898 857
rect 328 848 329 852
rect 331 848 332 852
rect 666 848 667 852
rect 669 848 670 852
rect 682 848 683 852
rect 685 848 686 852
rect 698 848 699 852
rect 701 848 702 852
rect 717 848 722 852
rect 724 848 727 852
rect 729 848 730 852
rect 751 848 753 852
rect 755 848 756 852
rect 773 848 774 852
rect 776 848 777 852
rect 789 848 794 852
rect 796 848 799 852
rect 801 848 802 852
rect 816 848 817 852
rect 819 848 820 852
rect 975 853 976 857
rect 978 853 979 857
rect 666 802 667 806
rect 669 802 670 806
rect 682 802 683 806
rect 685 802 686 806
rect 698 802 699 806
rect 701 802 702 806
rect 717 802 722 806
rect 724 802 727 806
rect 729 802 730 806
rect 751 802 753 806
rect 755 802 756 806
rect 773 802 774 806
rect 776 802 777 806
rect 789 802 794 806
rect 796 802 799 806
rect 801 802 802 806
rect 816 802 817 806
rect 819 802 820 806
rect 312 792 313 796
rect 315 792 316 796
rect 328 792 329 796
rect 331 792 334 796
rect 336 792 337 796
rect 349 792 350 796
rect 352 792 353 796
rect 365 792 366 796
rect 368 792 369 796
rect 386 792 387 796
rect 389 792 392 796
rect 394 792 395 796
rect 407 792 408 796
rect 410 792 411 796
rect 423 792 424 796
rect 426 792 429 796
rect 431 792 432 796
rect 864 801 867 805
rect 869 801 872 805
rect 874 801 875 805
rect 945 801 948 805
rect 950 801 953 805
rect 955 801 956 805
rect 864 725 867 729
rect 869 725 872 729
rect 874 725 875 729
rect 945 729 946 733
rect 948 729 949 733
rect 969 725 972 729
rect 974 725 977 729
rect 979 725 980 729
rect 894 721 895 725
rect 897 721 898 725
rect 666 716 667 720
rect 669 716 670 720
rect 682 716 683 720
rect 685 716 686 720
rect 698 716 699 720
rect 701 716 702 720
rect 717 716 722 720
rect 724 716 727 720
rect 729 716 730 720
rect 751 716 753 720
rect 755 716 756 720
rect 773 716 774 720
rect 776 716 777 720
rect 789 716 794 720
rect 796 716 799 720
rect 801 716 802 720
rect 816 716 817 720
rect 819 716 820 720
rect 999 721 1000 725
rect 1002 721 1003 725
rect 666 670 667 674
rect 669 670 670 674
rect 682 670 683 674
rect 685 670 686 674
rect 698 670 699 674
rect 701 670 702 674
rect 717 670 722 674
rect 724 670 727 674
rect 729 670 730 674
rect 751 670 753 674
rect 755 670 756 674
rect 773 670 774 674
rect 776 670 777 674
rect 789 670 794 674
rect 796 670 799 674
rect 801 670 802 674
rect 816 670 817 674
rect 819 670 820 674
rect 864 670 867 674
rect 869 670 872 674
rect 874 670 875 674
rect 969 670 972 674
rect 974 670 977 674
rect 979 670 980 674
rect 864 593 867 597
rect 869 593 872 597
rect 874 593 875 597
rect 921 597 922 601
rect 924 597 925 601
rect 945 593 948 597
rect 950 593 953 597
rect 955 593 956 597
rect 1011 597 1012 601
rect 1014 597 1015 601
rect 1035 593 1038 597
rect 1040 593 1043 597
rect 1045 593 1046 597
rect 894 589 895 593
rect 897 589 898 593
rect 666 584 667 588
rect 669 584 670 588
rect 682 584 683 588
rect 685 584 686 588
rect 698 584 699 588
rect 701 584 702 588
rect 717 584 722 588
rect 724 584 727 588
rect 729 584 730 588
rect 751 584 753 588
rect 755 584 756 588
rect 773 584 774 588
rect 776 584 777 588
rect 789 584 794 588
rect 796 584 799 588
rect 801 584 802 588
rect 816 584 817 588
rect 819 584 820 588
rect 975 589 976 593
rect 978 589 979 593
rect 1065 589 1066 593
rect 1068 589 1069 593
rect 666 538 667 542
rect 669 538 670 542
rect 682 538 683 542
rect 685 538 686 542
rect 698 538 699 542
rect 701 538 702 542
rect 717 538 722 542
rect 724 538 727 542
rect 729 538 730 542
rect 751 538 753 542
rect 755 538 756 542
rect 773 538 774 542
rect 776 538 777 542
rect 789 538 794 542
rect 796 538 799 542
rect 801 538 802 542
rect 816 538 817 542
rect 819 538 820 542
rect 864 535 867 539
rect 869 535 872 539
rect 874 535 875 539
rect 945 535 948 539
rect 950 535 953 539
rect 955 535 956 539
rect 1035 535 1038 539
rect 1040 535 1043 539
rect 1045 535 1046 539
rect 864 461 867 465
rect 869 461 872 465
rect 874 461 875 465
rect 894 457 895 461
rect 897 457 898 461
rect 666 452 667 456
rect 669 452 670 456
rect 682 452 683 456
rect 685 452 686 456
rect 698 452 699 456
rect 701 452 702 456
rect 717 452 722 456
rect 724 452 727 456
rect 729 452 730 456
rect 751 452 753 456
rect 755 452 756 456
rect 773 452 774 456
rect 776 452 777 456
rect 789 452 794 456
rect 796 452 799 456
rect 801 452 802 456
rect 816 452 817 456
rect 819 452 820 456
rect 666 406 667 410
rect 669 406 670 410
rect 682 406 683 410
rect 685 406 686 410
rect 698 406 699 410
rect 701 406 702 410
rect 717 406 722 410
rect 724 406 727 410
rect 729 406 730 410
rect 751 406 753 410
rect 755 406 756 410
rect 773 406 774 410
rect 776 406 777 410
rect 789 406 794 410
rect 796 406 799 410
rect 801 406 802 410
rect 816 406 817 410
rect 819 406 820 410
rect 900 406 901 410
rect 903 406 904 410
rect 908 406 914 410
rect 918 406 919 410
rect 921 406 922 410
rect 943 406 944 410
rect 946 406 947 410
rect 959 406 960 410
rect 962 406 963 410
rect 978 406 983 410
rect 985 406 988 410
rect 990 406 991 410
rect 1012 406 1014 410
rect 1016 406 1017 410
rect 1034 406 1035 410
rect 1037 406 1038 410
rect 1050 406 1055 410
rect 1057 406 1060 410
rect 1062 406 1063 410
rect 1077 406 1078 410
rect 1080 406 1081 410
rect 189 392 190 396
rect 192 392 195 396
rect 197 392 198 396
rect 210 392 211 396
rect 213 392 214 396
rect 226 392 227 396
rect 229 392 232 396
rect 234 392 235 396
rect 252 392 253 396
rect 255 392 256 396
rect 268 392 269 396
rect 271 392 272 396
rect 284 392 285 396
rect 287 392 290 396
rect 292 392 293 396
rect 305 392 306 396
rect 308 392 309 396
rect 321 392 322 396
rect 324 392 327 396
rect 329 392 330 396
rect 342 392 343 396
rect 345 392 346 396
rect 358 392 359 396
rect 361 392 364 396
rect 366 392 367 396
rect 384 392 385 396
rect 387 392 388 396
rect 400 392 401 396
rect 403 392 404 396
rect 416 392 417 396
rect 419 392 422 396
rect 424 392 425 396
rect 437 392 438 396
rect 440 392 441 396
rect 453 392 454 396
rect 456 392 459 396
rect 461 392 462 396
rect 474 392 475 396
rect 477 392 478 396
rect 490 392 491 396
rect 493 392 496 396
rect 498 392 499 396
rect 516 392 517 396
rect 519 392 520 396
rect 532 392 533 396
rect 535 392 536 396
rect 548 392 549 396
rect 551 392 554 396
rect 556 392 557 396
rect 569 392 570 396
rect 572 392 573 396
rect 864 399 867 403
rect 869 399 872 403
rect 874 399 875 403
rect 304 348 305 352
rect 307 348 308 352
rect 328 348 329 352
rect 331 348 332 352
rect 1090 352 1094 353
rect 1090 349 1094 350
rect 324 337 325 341
rect 327 337 328 341
rect 316 325 320 326
rect 316 322 320 323
rect 304 314 305 318
rect 307 314 308 318
rect 328 314 329 318
rect 331 314 332 318
rect 960 282 961 286
rect 963 282 966 286
rect 968 282 969 286
rect 981 282 982 286
rect 984 282 985 286
rect 997 282 998 286
rect 1000 282 1003 286
rect 1005 282 1006 286
rect 1023 282 1024 286
rect 1026 282 1027 286
rect 1039 282 1040 286
rect 1042 282 1043 286
rect 1055 282 1056 286
rect 1058 282 1061 286
rect 1063 282 1064 286
rect 1076 282 1077 286
rect 1079 282 1080 286
rect 189 252 190 256
rect 192 252 195 256
rect 197 252 198 256
rect 210 252 211 256
rect 213 252 214 256
rect 226 252 227 256
rect 229 252 232 256
rect 234 252 235 256
rect 252 252 253 256
rect 255 252 256 256
rect 268 252 269 256
rect 271 252 272 256
rect 284 252 285 256
rect 287 252 290 256
rect 292 252 293 256
rect 305 252 306 256
rect 308 252 309 256
rect 321 252 322 256
rect 324 252 327 256
rect 329 252 330 256
rect 342 252 343 256
rect 345 252 346 256
rect 358 252 359 256
rect 361 252 364 256
rect 366 252 367 256
rect 384 252 385 256
rect 387 252 388 256
rect 400 252 401 256
rect 403 252 404 256
rect 416 252 417 256
rect 419 252 422 256
rect 424 252 425 256
rect 437 252 438 256
rect 440 252 441 256
rect 453 252 454 256
rect 456 252 459 256
rect 461 252 462 256
rect 474 252 475 256
rect 477 252 478 256
rect 490 252 491 256
rect 493 252 496 256
rect 498 252 499 256
rect 516 252 517 256
rect 519 252 520 256
rect 532 252 533 256
rect 535 252 536 256
rect 548 252 549 256
rect 551 252 554 256
rect 556 252 557 256
rect 569 252 570 256
rect 572 252 573 256
rect 1102 208 1106 209
rect 1102 205 1106 206
rect 960 196 961 200
rect 963 196 966 200
rect 968 196 969 200
rect 981 196 982 200
rect 984 196 985 200
rect 997 196 998 200
rect 1000 196 1003 200
rect 1005 196 1006 200
rect 1023 196 1024 200
rect 1026 196 1027 200
rect 1039 196 1040 200
rect 1042 196 1043 200
rect 1055 196 1056 200
rect 1058 196 1061 200
rect 1063 196 1064 200
rect 1076 196 1077 200
rect 1079 196 1080 200
rect 189 166 190 170
rect 192 166 195 170
rect 197 166 198 170
rect 210 166 211 170
rect 213 166 214 170
rect 226 166 227 170
rect 229 166 232 170
rect 234 166 235 170
rect 252 166 253 170
rect 255 166 256 170
rect 268 166 269 170
rect 271 166 272 170
rect 284 166 285 170
rect 287 166 290 170
rect 292 166 293 170
rect 305 166 306 170
rect 308 166 309 170
rect 321 166 322 170
rect 324 166 327 170
rect 329 166 330 170
rect 342 166 343 170
rect 345 166 346 170
rect 358 166 359 170
rect 361 166 364 170
rect 366 166 367 170
rect 384 166 385 170
rect 387 166 388 170
rect 400 166 401 170
rect 403 166 404 170
rect 416 166 417 170
rect 419 166 422 170
rect 424 166 425 170
rect 437 166 438 170
rect 440 166 441 170
rect 453 166 454 170
rect 456 166 459 170
rect 461 166 462 170
rect 474 166 475 170
rect 477 166 478 170
rect 490 166 491 170
rect 493 166 496 170
rect 498 166 499 170
rect 516 166 517 170
rect 519 166 520 170
rect 532 166 533 170
rect 535 166 536 170
rect 548 166 549 170
rect 551 166 554 170
rect 556 166 557 170
rect 569 166 570 170
rect 572 166 573 170
rect 421 122 422 126
rect 424 122 425 126
rect 445 122 446 126
rect 448 122 449 126
rect 441 111 442 115
rect 444 111 445 115
rect 433 99 437 100
rect 433 96 437 97
rect 421 88 422 92
rect 424 88 425 92
rect 445 88 446 92
rect 448 88 449 92
rect 189 26 190 30
rect 192 26 195 30
rect 197 26 198 30
rect 210 26 211 30
rect 213 26 214 30
rect 226 26 227 30
rect 229 26 232 30
rect 234 26 235 30
rect 252 26 253 30
rect 255 26 256 30
rect 268 26 269 30
rect 271 26 272 30
rect 284 26 285 30
rect 287 26 290 30
rect 292 26 293 30
rect 305 26 306 30
rect 308 26 309 30
rect 321 26 322 30
rect 324 26 327 30
rect 329 26 330 30
rect 342 26 343 30
rect 345 26 346 30
rect 358 26 359 30
rect 361 26 364 30
rect 366 26 367 30
rect 384 26 385 30
rect 387 26 388 30
rect 400 26 401 30
rect 403 26 404 30
rect 416 26 417 30
rect 419 26 422 30
rect 424 26 425 30
rect 437 26 438 30
rect 440 26 441 30
rect 453 26 454 30
rect 456 26 459 30
rect 461 26 462 30
rect 474 26 475 30
rect 477 26 478 30
rect 490 26 491 30
rect 493 26 496 30
rect 498 26 499 30
rect 516 26 517 30
rect 519 26 520 30
rect 532 26 533 30
rect 535 26 536 30
rect 548 26 549 30
rect 551 26 554 30
rect 556 26 557 30
rect 569 26 570 30
rect 572 26 573 30
<< pdiffusion >>
rect 661 950 662 958
rect 664 950 667 958
rect 669 950 670 958
rect 682 950 683 958
rect 685 954 686 958
rect 685 950 690 954
rect 698 950 699 958
rect 701 950 704 958
rect 706 950 707 958
rect 724 950 725 958
rect 727 950 728 958
rect 740 950 741 958
rect 743 954 744 958
rect 743 950 748 954
rect 756 950 757 958
rect 759 950 762 958
rect 764 950 765 958
rect 777 950 778 958
rect 780 950 781 958
rect 793 950 794 958
rect 796 950 799 958
rect 801 950 802 958
rect 814 950 815 958
rect 817 954 818 958
rect 817 950 822 954
rect 830 950 831 958
rect 833 950 836 958
rect 838 950 839 958
rect 856 950 857 958
rect 859 950 860 958
rect 872 950 873 958
rect 875 954 876 958
rect 875 950 880 954
rect 888 950 889 958
rect 891 950 894 958
rect 896 950 897 958
rect 909 950 910 958
rect 912 950 913 958
rect 925 950 926 958
rect 928 950 931 958
rect 933 950 934 958
rect 946 950 947 958
rect 949 954 950 958
rect 949 950 954 954
rect 962 950 963 958
rect 965 950 968 958
rect 970 950 971 958
rect 988 950 989 958
rect 991 950 992 958
rect 1004 950 1005 958
rect 1007 954 1008 958
rect 1007 950 1012 954
rect 1020 950 1021 958
rect 1023 950 1026 958
rect 1028 950 1029 958
rect 1041 950 1042 958
rect 1044 950 1045 958
rect 1057 950 1058 958
rect 1060 950 1063 958
rect 1065 950 1066 958
rect 1078 950 1079 958
rect 1081 954 1082 958
rect 1081 950 1086 954
rect 1094 950 1095 958
rect 1097 950 1100 958
rect 1102 950 1103 958
rect 1120 950 1121 958
rect 1123 950 1124 958
rect 1136 950 1137 958
rect 1139 954 1140 958
rect 1139 950 1144 954
rect 1152 950 1153 958
rect 1155 950 1158 958
rect 1160 950 1161 958
rect 1173 950 1174 958
rect 1176 950 1177 958
rect 321 917 322 925
rect 324 917 327 925
rect 329 917 330 925
rect 342 917 343 925
rect 345 921 346 925
rect 345 917 350 921
rect 358 917 359 925
rect 361 917 364 925
rect 366 917 367 925
rect 384 917 385 925
rect 387 917 388 925
rect 400 917 401 925
rect 403 921 404 925
rect 403 917 408 921
rect 416 917 417 925
rect 419 917 422 925
rect 424 917 425 925
rect 437 917 438 925
rect 440 917 441 925
rect 840 879 841 887
rect 843 879 844 887
rect 666 866 667 874
rect 669 866 670 874
rect 682 866 683 874
rect 685 866 686 874
rect 698 866 699 874
rect 701 866 702 874
rect 717 866 722 874
rect 724 866 727 874
rect 729 866 730 874
rect 751 866 753 874
rect 755 866 756 874
rect 773 866 774 874
rect 776 866 777 874
rect 789 866 794 874
rect 796 866 799 874
rect 801 866 802 874
rect 816 866 817 874
rect 819 866 820 874
rect 864 873 867 881
rect 869 873 872 881
rect 874 873 875 881
rect 894 879 895 887
rect 897 879 898 887
rect 921 879 922 887
rect 924 879 925 887
rect 945 873 948 881
rect 950 873 953 881
rect 955 873 956 881
rect 975 879 976 887
rect 978 879 979 887
rect 312 815 313 823
rect 315 815 316 823
rect 328 815 329 823
rect 331 815 334 823
rect 336 815 337 823
rect 349 819 350 823
rect 345 815 350 819
rect 352 815 353 823
rect 365 815 366 823
rect 368 815 369 823
rect 386 815 387 823
rect 389 815 392 823
rect 394 815 395 823
rect 407 819 408 823
rect 403 815 408 819
rect 410 815 411 823
rect 423 815 424 823
rect 426 815 429 823
rect 431 815 432 823
rect 666 780 667 788
rect 669 780 670 788
rect 682 780 683 788
rect 685 780 686 788
rect 698 780 699 788
rect 701 780 702 788
rect 717 780 722 788
rect 724 780 727 788
rect 729 780 730 788
rect 751 780 753 788
rect 755 780 756 788
rect 773 780 774 788
rect 776 780 777 788
rect 789 780 794 788
rect 796 780 799 788
rect 801 780 802 788
rect 816 780 817 788
rect 819 780 820 788
rect 864 781 867 789
rect 869 781 872 789
rect 874 781 875 789
rect 945 781 948 789
rect 950 781 953 789
rect 955 781 956 789
rect 666 734 667 742
rect 669 734 670 742
rect 682 734 683 742
rect 685 734 686 742
rect 698 734 699 742
rect 701 734 702 742
rect 717 734 722 742
rect 724 734 727 742
rect 729 734 730 742
rect 751 734 753 742
rect 755 734 756 742
rect 773 734 774 742
rect 776 734 777 742
rect 789 734 794 742
rect 796 734 799 742
rect 801 734 802 742
rect 816 734 817 742
rect 819 734 820 742
rect 864 741 867 749
rect 869 741 872 749
rect 874 741 875 749
rect 894 747 895 755
rect 897 747 898 755
rect 945 747 946 755
rect 948 747 949 755
rect 969 741 972 749
rect 974 741 977 749
rect 979 741 980 749
rect 999 747 1000 755
rect 1002 747 1003 755
rect 666 648 667 656
rect 669 648 670 656
rect 682 648 683 656
rect 685 648 686 656
rect 698 648 699 656
rect 701 648 702 656
rect 717 648 722 656
rect 724 648 727 656
rect 729 648 730 656
rect 751 648 753 656
rect 755 648 756 656
rect 773 648 774 656
rect 776 648 777 656
rect 789 648 794 656
rect 796 648 799 656
rect 801 648 802 656
rect 816 648 817 656
rect 819 648 820 656
rect 864 650 867 658
rect 869 650 872 658
rect 874 650 875 658
rect 969 650 972 658
rect 974 650 977 658
rect 979 650 980 658
rect 666 602 667 610
rect 669 602 670 610
rect 682 602 683 610
rect 685 602 686 610
rect 698 602 699 610
rect 701 602 702 610
rect 717 602 722 610
rect 724 602 727 610
rect 729 602 730 610
rect 751 602 753 610
rect 755 602 756 610
rect 773 602 774 610
rect 776 602 777 610
rect 789 602 794 610
rect 796 602 799 610
rect 801 602 802 610
rect 816 602 817 610
rect 819 602 820 610
rect 864 609 867 617
rect 869 609 872 617
rect 874 609 875 617
rect 894 615 895 623
rect 897 615 898 623
rect 921 615 922 623
rect 924 615 925 623
rect 945 609 948 617
rect 950 609 953 617
rect 955 609 956 617
rect 975 615 976 623
rect 978 615 979 623
rect 1011 615 1012 623
rect 1014 615 1015 623
rect 1035 609 1038 617
rect 1040 609 1043 617
rect 1045 609 1046 617
rect 1065 615 1066 623
rect 1068 615 1069 623
rect 666 516 667 524
rect 669 516 670 524
rect 682 516 683 524
rect 685 516 686 524
rect 698 516 699 524
rect 701 516 702 524
rect 717 516 722 524
rect 724 516 727 524
rect 729 516 730 524
rect 751 516 753 524
rect 755 516 756 524
rect 773 516 774 524
rect 776 516 777 524
rect 789 516 794 524
rect 796 516 799 524
rect 801 516 802 524
rect 816 516 817 524
rect 819 516 820 524
rect 864 515 867 523
rect 869 515 872 523
rect 874 515 875 523
rect 945 515 948 523
rect 950 515 953 523
rect 955 515 956 523
rect 1035 515 1038 523
rect 1040 515 1043 523
rect 1045 515 1046 523
rect 666 470 667 478
rect 669 470 670 478
rect 682 470 683 478
rect 685 470 686 478
rect 698 470 699 478
rect 701 470 702 478
rect 717 470 722 478
rect 724 470 727 478
rect 729 470 730 478
rect 751 470 753 478
rect 755 470 756 478
rect 773 470 774 478
rect 776 470 777 478
rect 789 470 794 478
rect 796 470 799 478
rect 801 470 802 478
rect 816 470 817 478
rect 819 470 820 478
rect 864 477 867 485
rect 869 477 872 485
rect 874 477 875 485
rect 894 483 895 491
rect 897 483 898 491
rect 189 415 190 423
rect 192 415 195 423
rect 197 415 198 423
rect 210 415 211 423
rect 213 419 214 423
rect 213 415 218 419
rect 226 415 227 423
rect 229 415 232 423
rect 234 415 235 423
rect 252 415 253 423
rect 255 415 256 423
rect 268 415 269 423
rect 271 419 272 423
rect 271 415 276 419
rect 284 415 285 423
rect 287 415 290 423
rect 292 415 293 423
rect 305 415 306 423
rect 308 415 309 423
rect 321 415 322 423
rect 324 415 327 423
rect 329 415 330 423
rect 342 415 343 423
rect 345 419 346 423
rect 345 415 350 419
rect 358 415 359 423
rect 361 415 364 423
rect 366 415 367 423
rect 384 415 385 423
rect 387 415 388 423
rect 400 415 401 423
rect 403 419 404 423
rect 403 415 408 419
rect 416 415 417 423
rect 419 415 422 423
rect 424 415 425 423
rect 437 415 438 423
rect 440 415 441 423
rect 453 415 454 423
rect 456 415 459 423
rect 461 415 462 423
rect 474 415 475 423
rect 477 419 478 423
rect 477 415 482 419
rect 490 415 491 423
rect 493 415 496 423
rect 498 415 499 423
rect 516 415 517 423
rect 519 415 520 423
rect 532 415 533 423
rect 535 419 536 423
rect 535 415 540 419
rect 548 415 549 423
rect 551 415 554 423
rect 556 415 557 423
rect 569 415 570 423
rect 572 415 573 423
rect 666 384 667 392
rect 669 384 670 392
rect 682 384 683 392
rect 685 384 686 392
rect 698 384 699 392
rect 701 384 702 392
rect 717 384 722 392
rect 724 384 727 392
rect 729 384 730 392
rect 751 384 753 392
rect 755 384 756 392
rect 773 384 774 392
rect 776 384 777 392
rect 789 384 794 392
rect 796 384 799 392
rect 801 384 802 392
rect 816 384 817 392
rect 819 384 820 392
rect 864 379 867 387
rect 869 379 872 387
rect 874 379 875 387
rect 900 384 901 392
rect 903 384 904 392
rect 908 384 914 392
rect 918 384 919 392
rect 921 384 922 392
rect 943 384 944 392
rect 946 384 947 392
rect 959 384 960 392
rect 962 384 963 392
rect 978 384 983 392
rect 985 384 988 392
rect 990 384 991 392
rect 1012 384 1014 392
rect 1016 384 1017 392
rect 1034 384 1035 392
rect 1037 384 1038 392
rect 1050 384 1055 392
rect 1057 384 1060 392
rect 1062 384 1063 392
rect 1077 384 1078 392
rect 1080 384 1081 392
rect 960 305 961 313
rect 963 305 966 313
rect 968 305 969 313
rect 981 305 982 313
rect 984 309 985 313
rect 984 305 989 309
rect 997 305 998 313
rect 1000 305 1003 313
rect 1005 305 1006 313
rect 1023 305 1024 313
rect 1026 305 1027 313
rect 1039 305 1040 313
rect 1042 309 1043 313
rect 1042 305 1047 309
rect 1055 305 1056 313
rect 1058 305 1061 313
rect 1063 305 1064 313
rect 1076 305 1077 313
rect 1079 305 1080 313
rect 189 275 190 283
rect 192 275 195 283
rect 197 275 198 283
rect 210 275 211 283
rect 213 279 214 283
rect 213 275 218 279
rect 226 275 227 283
rect 229 275 232 283
rect 234 275 235 283
rect 252 275 253 283
rect 255 275 256 283
rect 268 275 269 283
rect 271 279 272 283
rect 271 275 276 279
rect 284 275 285 283
rect 287 275 290 283
rect 292 275 293 283
rect 305 275 306 283
rect 308 275 309 283
rect 321 275 322 283
rect 324 275 327 283
rect 329 275 330 283
rect 342 275 343 283
rect 345 279 346 283
rect 345 275 350 279
rect 358 275 359 283
rect 361 275 364 283
rect 366 275 367 283
rect 384 275 385 283
rect 387 275 388 283
rect 400 275 401 283
rect 403 279 404 283
rect 403 275 408 279
rect 416 275 417 283
rect 419 275 422 283
rect 424 275 425 283
rect 437 275 438 283
rect 440 275 441 283
rect 453 275 454 283
rect 456 275 459 283
rect 461 275 462 283
rect 474 275 475 283
rect 477 279 478 283
rect 477 275 482 279
rect 490 275 491 283
rect 493 275 496 283
rect 498 275 499 283
rect 516 275 517 283
rect 519 275 520 283
rect 532 275 533 283
rect 535 279 536 283
rect 535 275 540 279
rect 548 275 549 283
rect 551 275 554 283
rect 556 275 557 283
rect 569 275 570 283
rect 572 275 573 283
rect 960 219 961 227
rect 963 219 966 227
rect 968 219 969 227
rect 981 219 982 227
rect 984 223 985 227
rect 984 219 989 223
rect 997 219 998 227
rect 1000 219 1003 227
rect 1005 219 1006 227
rect 1023 219 1024 227
rect 1026 219 1027 227
rect 1039 219 1040 227
rect 1042 223 1043 227
rect 1042 219 1047 223
rect 1055 219 1056 227
rect 1058 219 1061 227
rect 1063 219 1064 227
rect 1076 219 1077 227
rect 1079 219 1080 227
rect 189 189 190 197
rect 192 189 195 197
rect 197 189 198 197
rect 210 189 211 197
rect 213 193 214 197
rect 213 189 218 193
rect 226 189 227 197
rect 229 189 232 197
rect 234 189 235 197
rect 252 189 253 197
rect 255 189 256 197
rect 268 189 269 197
rect 271 193 272 197
rect 271 189 276 193
rect 284 189 285 197
rect 287 189 290 197
rect 292 189 293 197
rect 305 189 306 197
rect 308 189 309 197
rect 321 189 322 197
rect 324 189 327 197
rect 329 189 330 197
rect 342 189 343 197
rect 345 193 346 197
rect 345 189 350 193
rect 358 189 359 197
rect 361 189 364 197
rect 366 189 367 197
rect 384 189 385 197
rect 387 189 388 197
rect 400 189 401 197
rect 403 193 404 197
rect 403 189 408 193
rect 416 189 417 197
rect 419 189 422 197
rect 424 189 425 197
rect 437 189 438 197
rect 440 189 441 197
rect 453 189 454 197
rect 456 189 459 197
rect 461 189 462 197
rect 474 189 475 197
rect 477 193 478 197
rect 477 189 482 193
rect 490 189 491 197
rect 493 189 496 197
rect 498 189 499 197
rect 516 189 517 197
rect 519 189 520 197
rect 532 189 533 197
rect 535 193 536 197
rect 535 189 540 193
rect 548 189 549 197
rect 551 189 554 197
rect 556 189 557 197
rect 569 189 570 197
rect 572 189 573 197
rect 189 49 190 57
rect 192 49 195 57
rect 197 49 198 57
rect 210 49 211 57
rect 213 53 214 57
rect 213 49 218 53
rect 226 49 227 57
rect 229 49 232 57
rect 234 49 235 57
rect 252 49 253 57
rect 255 49 256 57
rect 268 49 269 57
rect 271 53 272 57
rect 271 49 276 53
rect 284 49 285 57
rect 287 49 290 57
rect 292 49 293 57
rect 305 49 306 57
rect 308 49 309 57
rect 321 49 322 57
rect 324 49 327 57
rect 329 49 330 57
rect 342 49 343 57
rect 345 53 346 57
rect 345 49 350 53
rect 358 49 359 57
rect 361 49 364 57
rect 366 49 367 57
rect 384 49 385 57
rect 387 49 388 57
rect 400 49 401 57
rect 403 53 404 57
rect 403 49 408 53
rect 416 49 417 57
rect 419 49 422 57
rect 424 49 425 57
rect 437 49 438 57
rect 440 49 441 57
rect 453 49 454 57
rect 456 49 459 57
rect 461 49 462 57
rect 474 49 475 57
rect 477 53 478 57
rect 477 49 482 53
rect 490 49 491 57
rect 493 49 496 57
rect 498 49 499 57
rect 516 49 517 57
rect 519 49 520 57
rect 532 49 533 57
rect 535 53 536 57
rect 535 49 540 53
rect 548 49 549 57
rect 551 49 554 57
rect 556 49 557 57
rect 569 49 570 57
rect 572 49 573 57
<< ndcontact >>
rect 657 927 661 931
rect 670 927 674 931
rect 678 927 682 931
rect 686 927 690 931
rect 694 927 698 931
rect 707 927 711 931
rect 720 927 724 931
rect 728 927 732 931
rect 736 927 740 931
rect 744 927 748 931
rect 752 927 756 931
rect 765 927 769 931
rect 773 927 777 931
rect 781 927 785 931
rect 789 927 793 931
rect 802 927 806 931
rect 810 927 814 931
rect 818 927 822 931
rect 826 927 830 931
rect 839 927 843 931
rect 852 927 856 931
rect 860 927 864 931
rect 868 927 872 931
rect 876 927 880 931
rect 884 927 888 931
rect 897 927 901 931
rect 905 927 909 931
rect 913 927 917 931
rect 921 927 925 931
rect 934 927 938 931
rect 942 927 946 931
rect 950 927 954 931
rect 958 927 962 931
rect 971 927 975 931
rect 984 927 988 931
rect 992 927 996 931
rect 1000 927 1004 931
rect 1008 927 1012 931
rect 1016 927 1020 931
rect 1029 927 1033 931
rect 1037 927 1041 931
rect 1045 927 1049 931
rect 1053 927 1057 931
rect 1066 927 1070 931
rect 1074 927 1078 931
rect 1082 927 1086 931
rect 1090 927 1094 931
rect 1103 927 1107 931
rect 1116 927 1120 931
rect 1124 927 1128 931
rect 1132 927 1136 931
rect 1140 927 1144 931
rect 1148 927 1152 931
rect 1161 927 1165 931
rect 1169 927 1173 931
rect 1177 927 1181 931
rect 317 894 321 898
rect 330 894 334 898
rect 338 894 342 898
rect 346 894 350 898
rect 354 894 358 898
rect 367 894 371 898
rect 380 894 384 898
rect 388 894 392 898
rect 396 894 400 898
rect 404 894 408 898
rect 412 894 416 898
rect 425 894 429 898
rect 433 894 437 898
rect 441 894 445 898
rect 441 857 445 861
rect 449 857 453 861
rect 836 861 840 865
rect 844 861 848 865
rect 860 857 864 861
rect 875 857 879 861
rect 917 861 921 865
rect 925 861 929 865
rect 941 857 945 861
rect 956 857 960 861
rect 890 853 894 857
rect 898 853 902 857
rect 324 848 328 852
rect 332 848 336 852
rect 662 848 666 852
rect 670 848 674 852
rect 678 848 682 852
rect 686 848 690 852
rect 694 848 698 852
rect 702 848 706 852
rect 713 848 717 852
rect 730 848 734 852
rect 747 848 751 852
rect 756 848 760 852
rect 769 848 773 852
rect 777 848 781 852
rect 785 848 789 852
rect 802 848 806 852
rect 812 848 816 852
rect 820 848 824 852
rect 971 853 975 857
rect 979 853 983 857
rect 662 802 666 806
rect 670 802 674 806
rect 678 802 682 806
rect 686 802 690 806
rect 694 802 698 806
rect 702 802 706 806
rect 713 802 717 806
rect 730 802 734 806
rect 747 802 751 806
rect 756 802 760 806
rect 769 802 773 806
rect 777 802 781 806
rect 785 802 789 806
rect 802 802 806 806
rect 812 802 816 806
rect 820 802 824 806
rect 308 792 312 796
rect 316 792 320 796
rect 324 792 328 796
rect 337 792 341 796
rect 345 792 349 796
rect 353 792 357 796
rect 361 792 365 796
rect 369 792 373 796
rect 382 792 386 796
rect 395 792 399 796
rect 403 792 407 796
rect 411 792 415 796
rect 419 792 423 796
rect 432 792 436 796
rect 860 801 864 805
rect 875 801 879 805
rect 941 801 945 805
rect 956 801 960 805
rect 860 725 864 729
rect 875 725 879 729
rect 941 729 945 733
rect 949 729 953 733
rect 965 725 969 729
rect 980 725 984 729
rect 890 721 894 725
rect 898 721 902 725
rect 662 716 666 720
rect 670 716 674 720
rect 678 716 682 720
rect 686 716 690 720
rect 694 716 698 720
rect 702 716 706 720
rect 713 716 717 720
rect 730 716 734 720
rect 747 716 751 720
rect 756 716 760 720
rect 769 716 773 720
rect 777 716 781 720
rect 785 716 789 720
rect 802 716 806 720
rect 812 716 816 720
rect 820 716 824 720
rect 995 721 999 725
rect 1003 721 1007 725
rect 662 670 666 674
rect 670 670 674 674
rect 678 670 682 674
rect 686 670 690 674
rect 694 670 698 674
rect 702 670 706 674
rect 713 670 717 674
rect 730 670 734 674
rect 747 670 751 674
rect 756 670 760 674
rect 769 670 773 674
rect 777 670 781 674
rect 785 670 789 674
rect 802 670 806 674
rect 812 670 816 674
rect 820 670 824 674
rect 860 670 864 674
rect 875 670 879 674
rect 965 670 969 674
rect 980 670 984 674
rect 860 593 864 597
rect 875 593 879 597
rect 917 597 921 601
rect 925 597 929 601
rect 941 593 945 597
rect 956 593 960 597
rect 1007 597 1011 601
rect 1015 597 1019 601
rect 1031 593 1035 597
rect 1046 593 1050 597
rect 890 589 894 593
rect 898 589 902 593
rect 662 584 666 588
rect 670 584 674 588
rect 678 584 682 588
rect 686 584 690 588
rect 694 584 698 588
rect 702 584 706 588
rect 713 584 717 588
rect 730 584 734 588
rect 747 584 751 588
rect 756 584 760 588
rect 769 584 773 588
rect 777 584 781 588
rect 785 584 789 588
rect 802 584 806 588
rect 812 584 816 588
rect 820 584 824 588
rect 971 589 975 593
rect 979 589 983 593
rect 1061 589 1065 593
rect 1069 589 1073 593
rect 662 538 666 542
rect 670 538 674 542
rect 678 538 682 542
rect 686 538 690 542
rect 694 538 698 542
rect 702 538 706 542
rect 713 538 717 542
rect 730 538 734 542
rect 747 538 751 542
rect 756 538 760 542
rect 769 538 773 542
rect 777 538 781 542
rect 785 538 789 542
rect 802 538 806 542
rect 812 538 816 542
rect 820 538 824 542
rect 860 535 864 539
rect 875 535 879 539
rect 941 535 945 539
rect 956 535 960 539
rect 1031 535 1035 539
rect 1046 535 1050 539
rect 860 461 864 465
rect 875 461 879 465
rect 890 457 894 461
rect 898 457 902 461
rect 662 452 666 456
rect 670 452 674 456
rect 678 452 682 456
rect 686 452 690 456
rect 694 452 698 456
rect 702 452 706 456
rect 713 452 717 456
rect 730 452 734 456
rect 747 452 751 456
rect 756 452 760 456
rect 769 452 773 456
rect 777 452 781 456
rect 785 452 789 456
rect 802 452 806 456
rect 812 452 816 456
rect 820 452 824 456
rect 662 406 666 410
rect 670 406 674 410
rect 678 406 682 410
rect 686 406 690 410
rect 694 406 698 410
rect 702 406 706 410
rect 713 406 717 410
rect 730 406 734 410
rect 747 406 751 410
rect 756 406 760 410
rect 769 406 773 410
rect 777 406 781 410
rect 785 406 789 410
rect 802 406 806 410
rect 812 406 816 410
rect 820 406 824 410
rect 896 406 900 410
rect 904 406 908 410
rect 914 406 918 410
rect 922 406 926 410
rect 931 406 935 410
rect 939 406 943 410
rect 947 406 951 410
rect 955 406 959 410
rect 963 406 967 410
rect 974 406 978 410
rect 991 406 995 410
rect 1008 406 1012 410
rect 1017 406 1021 410
rect 1030 406 1034 410
rect 1038 406 1042 410
rect 1046 406 1050 410
rect 1063 406 1067 410
rect 1073 406 1077 410
rect 1081 406 1085 410
rect 185 392 189 396
rect 198 392 202 396
rect 206 392 210 396
rect 214 392 218 396
rect 222 392 226 396
rect 235 392 239 396
rect 248 392 252 396
rect 256 392 260 396
rect 264 392 268 396
rect 272 392 276 396
rect 280 392 284 396
rect 293 392 297 396
rect 301 392 305 396
rect 309 392 313 396
rect 317 392 321 396
rect 330 392 334 396
rect 338 392 342 396
rect 346 392 350 396
rect 354 392 358 396
rect 367 392 371 396
rect 380 392 384 396
rect 388 392 392 396
rect 396 392 400 396
rect 404 392 408 396
rect 412 392 416 396
rect 425 392 429 396
rect 433 392 437 396
rect 441 392 445 396
rect 449 392 453 396
rect 462 392 466 396
rect 470 392 474 396
rect 478 392 482 396
rect 486 392 490 396
rect 499 392 503 396
rect 512 392 516 396
rect 520 392 524 396
rect 528 392 532 396
rect 536 392 540 396
rect 544 392 548 396
rect 557 392 561 396
rect 565 392 569 396
rect 573 392 577 396
rect 860 399 864 403
rect 875 399 879 403
rect 1090 353 1094 357
rect 300 348 304 352
rect 308 348 312 352
rect 324 348 328 352
rect 332 348 336 352
rect 1090 345 1094 349
rect 320 337 324 341
rect 328 337 332 341
rect 316 326 320 330
rect 316 318 320 322
rect 300 314 304 318
rect 308 314 312 318
rect 324 314 328 318
rect 332 314 336 318
rect 956 282 960 286
rect 969 282 973 286
rect 977 282 981 286
rect 985 282 989 286
rect 993 282 997 286
rect 1006 282 1010 286
rect 1019 282 1023 286
rect 1027 282 1031 286
rect 1035 282 1039 286
rect 1043 282 1047 286
rect 1051 282 1055 286
rect 1064 282 1068 286
rect 1072 282 1076 286
rect 1080 282 1084 286
rect 185 252 189 256
rect 198 252 202 256
rect 206 252 210 256
rect 214 252 218 256
rect 222 252 226 256
rect 235 252 239 256
rect 248 252 252 256
rect 256 252 260 256
rect 264 252 268 256
rect 272 252 276 256
rect 280 252 284 256
rect 293 252 297 256
rect 301 252 305 256
rect 309 252 313 256
rect 317 252 321 256
rect 330 252 334 256
rect 338 252 342 256
rect 346 252 350 256
rect 354 252 358 256
rect 367 252 371 256
rect 380 252 384 256
rect 388 252 392 256
rect 396 252 400 256
rect 404 252 408 256
rect 412 252 416 256
rect 425 252 429 256
rect 433 252 437 256
rect 441 252 445 256
rect 449 252 453 256
rect 462 252 466 256
rect 470 252 474 256
rect 478 252 482 256
rect 486 252 490 256
rect 499 252 503 256
rect 512 252 516 256
rect 520 252 524 256
rect 528 252 532 256
rect 536 252 540 256
rect 544 252 548 256
rect 557 252 561 256
rect 565 252 569 256
rect 573 252 577 256
rect 1102 209 1106 213
rect 1102 201 1106 205
rect 956 196 960 200
rect 969 196 973 200
rect 977 196 981 200
rect 985 196 989 200
rect 993 196 997 200
rect 1006 196 1010 200
rect 1019 196 1023 200
rect 1027 196 1031 200
rect 1035 196 1039 200
rect 1043 196 1047 200
rect 1051 196 1055 200
rect 1064 196 1068 200
rect 1072 196 1076 200
rect 1080 196 1084 200
rect 185 166 189 170
rect 198 166 202 170
rect 206 166 210 170
rect 214 166 218 170
rect 222 166 226 170
rect 235 166 239 170
rect 248 166 252 170
rect 256 166 260 170
rect 264 166 268 170
rect 272 166 276 170
rect 280 166 284 170
rect 293 166 297 170
rect 301 166 305 170
rect 309 166 313 170
rect 317 166 321 170
rect 330 166 334 170
rect 338 166 342 170
rect 346 166 350 170
rect 354 166 358 170
rect 367 166 371 170
rect 380 166 384 170
rect 388 166 392 170
rect 396 166 400 170
rect 404 166 408 170
rect 412 166 416 170
rect 425 166 429 170
rect 433 166 437 170
rect 441 166 445 170
rect 449 166 453 170
rect 462 166 466 170
rect 470 166 474 170
rect 478 166 482 170
rect 486 166 490 170
rect 499 166 503 170
rect 512 166 516 170
rect 520 166 524 170
rect 528 166 532 170
rect 536 166 540 170
rect 544 166 548 170
rect 557 166 561 170
rect 565 166 569 170
rect 573 166 577 170
rect 417 122 421 126
rect 425 122 429 126
rect 441 122 445 126
rect 449 122 453 126
rect 437 111 441 115
rect 445 111 449 115
rect 433 100 437 104
rect 433 92 437 96
rect 417 88 421 92
rect 425 88 429 92
rect 441 88 445 92
rect 449 88 453 92
rect 185 26 189 30
rect 198 26 202 30
rect 206 26 210 30
rect 214 26 218 30
rect 222 26 226 30
rect 235 26 239 30
rect 248 26 252 30
rect 256 26 260 30
rect 264 26 268 30
rect 272 26 276 30
rect 280 26 284 30
rect 293 26 297 30
rect 301 26 305 30
rect 309 26 313 30
rect 317 26 321 30
rect 330 26 334 30
rect 338 26 342 30
rect 346 26 350 30
rect 354 26 358 30
rect 367 26 371 30
rect 380 26 384 30
rect 388 26 392 30
rect 396 26 400 30
rect 404 26 408 30
rect 412 26 416 30
rect 425 26 429 30
rect 433 26 437 30
rect 441 26 445 30
rect 449 26 453 30
rect 462 26 466 30
rect 470 26 474 30
rect 478 26 482 30
rect 486 26 490 30
rect 499 26 503 30
rect 512 26 516 30
rect 520 26 524 30
rect 528 26 532 30
rect 536 26 540 30
rect 544 26 548 30
rect 557 26 561 30
rect 565 26 569 30
rect 573 26 577 30
<< pdcontact >>
rect 657 950 661 958
rect 670 950 674 958
rect 678 950 682 958
rect 686 954 690 958
rect 694 950 698 958
rect 707 950 711 958
rect 720 950 724 958
rect 728 950 732 958
rect 736 950 740 958
rect 744 954 748 958
rect 752 950 756 958
rect 765 950 769 958
rect 773 950 777 958
rect 781 950 785 958
rect 789 950 793 958
rect 802 950 806 958
rect 810 950 814 958
rect 818 954 822 958
rect 826 950 830 958
rect 839 950 843 958
rect 852 950 856 958
rect 860 950 864 958
rect 868 950 872 958
rect 876 954 880 958
rect 884 950 888 958
rect 897 950 901 958
rect 905 950 909 958
rect 913 950 917 958
rect 921 950 925 958
rect 934 950 938 958
rect 942 950 946 958
rect 950 954 954 958
rect 958 950 962 958
rect 971 950 975 958
rect 984 950 988 958
rect 992 950 996 958
rect 1000 950 1004 958
rect 1008 954 1012 958
rect 1016 950 1020 958
rect 1029 950 1033 958
rect 1037 950 1041 958
rect 1045 950 1049 958
rect 1053 950 1057 958
rect 1066 950 1070 958
rect 1074 950 1078 958
rect 1082 954 1086 958
rect 1090 950 1094 958
rect 1103 950 1107 958
rect 1116 950 1120 958
rect 1124 950 1128 958
rect 1132 950 1136 958
rect 1140 954 1144 958
rect 1148 950 1152 958
rect 1161 950 1165 958
rect 1169 950 1173 958
rect 1177 950 1181 958
rect 317 917 321 925
rect 330 917 334 925
rect 338 917 342 925
rect 346 921 350 925
rect 354 917 358 925
rect 367 917 371 925
rect 380 917 384 925
rect 388 917 392 925
rect 396 917 400 925
rect 404 921 408 925
rect 412 917 416 925
rect 425 917 429 925
rect 433 917 437 925
rect 441 917 445 925
rect 836 879 840 887
rect 844 879 848 887
rect 662 866 666 874
rect 670 866 674 874
rect 678 866 682 874
rect 686 866 690 874
rect 694 866 698 874
rect 702 866 706 874
rect 713 866 717 874
rect 730 866 734 874
rect 747 866 751 874
rect 756 866 760 874
rect 769 866 773 874
rect 777 866 781 874
rect 785 866 789 874
rect 802 866 806 874
rect 812 866 816 874
rect 820 866 824 874
rect 860 873 864 881
rect 875 873 879 881
rect 890 879 894 887
rect 898 879 902 887
rect 917 879 921 887
rect 925 879 929 887
rect 941 873 945 881
rect 956 873 960 881
rect 971 879 975 887
rect 979 879 983 887
rect 308 815 312 823
rect 316 815 320 823
rect 324 815 328 823
rect 337 815 341 823
rect 345 819 349 823
rect 353 815 357 823
rect 361 815 365 823
rect 369 815 373 823
rect 382 815 386 823
rect 395 815 399 823
rect 403 819 407 823
rect 411 815 415 823
rect 419 815 423 823
rect 432 815 436 823
rect 662 780 666 788
rect 670 780 674 788
rect 678 780 682 788
rect 686 780 690 788
rect 694 780 698 788
rect 702 780 706 788
rect 713 780 717 788
rect 730 780 734 788
rect 747 780 751 788
rect 756 780 760 788
rect 769 780 773 788
rect 777 780 781 788
rect 785 780 789 788
rect 802 780 806 788
rect 812 780 816 788
rect 820 780 824 788
rect 860 781 864 789
rect 875 781 879 789
rect 941 781 945 789
rect 956 781 960 789
rect 662 734 666 742
rect 670 734 674 742
rect 678 734 682 742
rect 686 734 690 742
rect 694 734 698 742
rect 702 734 706 742
rect 713 734 717 742
rect 730 734 734 742
rect 747 734 751 742
rect 756 734 760 742
rect 769 734 773 742
rect 777 734 781 742
rect 785 734 789 742
rect 802 734 806 742
rect 812 734 816 742
rect 820 734 824 742
rect 860 741 864 749
rect 875 741 879 749
rect 890 747 894 755
rect 898 747 902 755
rect 941 747 945 755
rect 949 747 953 755
rect 965 741 969 749
rect 980 741 984 749
rect 995 747 999 755
rect 1003 747 1007 755
rect 662 648 666 656
rect 670 648 674 656
rect 678 648 682 656
rect 686 648 690 656
rect 694 648 698 656
rect 702 648 706 656
rect 713 648 717 656
rect 730 648 734 656
rect 747 648 751 656
rect 756 648 760 656
rect 769 648 773 656
rect 777 648 781 656
rect 785 648 789 656
rect 802 648 806 656
rect 812 648 816 656
rect 820 648 824 656
rect 860 650 864 658
rect 875 650 879 658
rect 965 650 969 658
rect 980 650 984 658
rect 662 602 666 610
rect 670 602 674 610
rect 678 602 682 610
rect 686 602 690 610
rect 694 602 698 610
rect 702 602 706 610
rect 713 602 717 610
rect 730 602 734 610
rect 747 602 751 610
rect 756 602 760 610
rect 769 602 773 610
rect 777 602 781 610
rect 785 602 789 610
rect 802 602 806 610
rect 812 602 816 610
rect 820 602 824 610
rect 860 609 864 617
rect 875 609 879 617
rect 890 615 894 623
rect 898 615 902 623
rect 917 615 921 623
rect 925 615 929 623
rect 941 609 945 617
rect 956 609 960 617
rect 971 615 975 623
rect 979 615 983 623
rect 1007 615 1011 623
rect 1015 615 1019 623
rect 1031 609 1035 617
rect 1046 609 1050 617
rect 1061 615 1065 623
rect 1069 615 1073 623
rect 662 516 666 524
rect 670 516 674 524
rect 678 516 682 524
rect 686 516 690 524
rect 694 516 698 524
rect 702 516 706 524
rect 713 516 717 524
rect 730 516 734 524
rect 747 516 751 524
rect 756 516 760 524
rect 769 516 773 524
rect 777 516 781 524
rect 785 516 789 524
rect 802 516 806 524
rect 812 516 816 524
rect 820 516 824 524
rect 860 515 864 523
rect 875 515 879 523
rect 941 515 945 523
rect 956 515 960 523
rect 1031 515 1035 523
rect 1046 515 1050 523
rect 662 470 666 478
rect 670 470 674 478
rect 678 470 682 478
rect 686 470 690 478
rect 694 470 698 478
rect 702 470 706 478
rect 713 470 717 478
rect 730 470 734 478
rect 747 470 751 478
rect 756 470 760 478
rect 769 470 773 478
rect 777 470 781 478
rect 785 470 789 478
rect 802 470 806 478
rect 812 470 816 478
rect 820 470 824 478
rect 860 477 864 485
rect 875 477 879 485
rect 890 483 894 491
rect 898 483 902 491
rect 185 415 189 423
rect 198 415 202 423
rect 206 415 210 423
rect 214 419 218 423
rect 222 415 226 423
rect 235 415 239 423
rect 248 415 252 423
rect 256 415 260 423
rect 264 415 268 423
rect 272 419 276 423
rect 280 415 284 423
rect 293 415 297 423
rect 301 415 305 423
rect 309 415 313 423
rect 317 415 321 423
rect 330 415 334 423
rect 338 415 342 423
rect 346 419 350 423
rect 354 415 358 423
rect 367 415 371 423
rect 380 415 384 423
rect 388 415 392 423
rect 396 415 400 423
rect 404 419 408 423
rect 412 415 416 423
rect 425 415 429 423
rect 433 415 437 423
rect 441 415 445 423
rect 449 415 453 423
rect 462 415 466 423
rect 470 415 474 423
rect 478 419 482 423
rect 486 415 490 423
rect 499 415 503 423
rect 512 415 516 423
rect 520 415 524 423
rect 528 415 532 423
rect 536 419 540 423
rect 544 415 548 423
rect 557 415 561 423
rect 565 415 569 423
rect 573 415 577 423
rect 662 384 666 392
rect 670 384 674 392
rect 678 384 682 392
rect 686 384 690 392
rect 694 384 698 392
rect 702 384 706 392
rect 713 384 717 392
rect 730 384 734 392
rect 747 384 751 392
rect 756 384 760 392
rect 769 384 773 392
rect 777 384 781 392
rect 785 384 789 392
rect 802 384 806 392
rect 812 384 816 392
rect 820 384 824 392
rect 860 379 864 387
rect 875 379 879 387
rect 896 384 900 392
rect 904 384 908 392
rect 914 384 918 392
rect 922 384 926 392
rect 931 384 935 392
rect 939 384 943 392
rect 947 384 951 392
rect 955 384 959 392
rect 963 384 967 392
rect 974 384 978 392
rect 991 384 995 392
rect 1008 384 1012 392
rect 1017 384 1021 392
rect 1030 384 1034 392
rect 1038 384 1042 392
rect 1046 384 1050 392
rect 1063 384 1067 392
rect 1073 384 1077 392
rect 1081 384 1085 392
rect 956 305 960 313
rect 969 305 973 313
rect 977 305 981 313
rect 985 309 989 313
rect 993 305 997 313
rect 1006 305 1010 313
rect 1019 305 1023 313
rect 1027 305 1031 313
rect 1035 305 1039 313
rect 1043 309 1047 313
rect 1051 305 1055 313
rect 1064 305 1068 313
rect 1072 305 1076 313
rect 1080 305 1084 313
rect 185 275 189 283
rect 198 275 202 283
rect 206 275 210 283
rect 214 279 218 283
rect 222 275 226 283
rect 235 275 239 283
rect 248 275 252 283
rect 256 275 260 283
rect 264 275 268 283
rect 272 279 276 283
rect 280 275 284 283
rect 293 275 297 283
rect 301 275 305 283
rect 309 275 313 283
rect 317 275 321 283
rect 330 275 334 283
rect 338 275 342 283
rect 346 279 350 283
rect 354 275 358 283
rect 367 275 371 283
rect 380 275 384 283
rect 388 275 392 283
rect 396 275 400 283
rect 404 279 408 283
rect 412 275 416 283
rect 425 275 429 283
rect 433 275 437 283
rect 441 275 445 283
rect 449 275 453 283
rect 462 275 466 283
rect 470 275 474 283
rect 478 279 482 283
rect 486 275 490 283
rect 499 275 503 283
rect 512 275 516 283
rect 520 275 524 283
rect 528 275 532 283
rect 536 279 540 283
rect 544 275 548 283
rect 557 275 561 283
rect 565 275 569 283
rect 573 275 577 283
rect 956 219 960 227
rect 969 219 973 227
rect 977 219 981 227
rect 985 223 989 227
rect 993 219 997 227
rect 1006 219 1010 227
rect 1019 219 1023 227
rect 1027 219 1031 227
rect 1035 219 1039 227
rect 1043 223 1047 227
rect 1051 219 1055 227
rect 1064 219 1068 227
rect 1072 219 1076 227
rect 1080 219 1084 227
rect 185 189 189 197
rect 198 189 202 197
rect 206 189 210 197
rect 214 193 218 197
rect 222 189 226 197
rect 235 189 239 197
rect 248 189 252 197
rect 256 189 260 197
rect 264 189 268 197
rect 272 193 276 197
rect 280 189 284 197
rect 293 189 297 197
rect 301 189 305 197
rect 309 189 313 197
rect 317 189 321 197
rect 330 189 334 197
rect 338 189 342 197
rect 346 193 350 197
rect 354 189 358 197
rect 367 189 371 197
rect 380 189 384 197
rect 388 189 392 197
rect 396 189 400 197
rect 404 193 408 197
rect 412 189 416 197
rect 425 189 429 197
rect 433 189 437 197
rect 441 189 445 197
rect 449 189 453 197
rect 462 189 466 197
rect 470 189 474 197
rect 478 193 482 197
rect 486 189 490 197
rect 499 189 503 197
rect 512 189 516 197
rect 520 189 524 197
rect 528 189 532 197
rect 536 193 540 197
rect 544 189 548 197
rect 557 189 561 197
rect 565 189 569 197
rect 573 189 577 197
rect 185 49 189 57
rect 198 49 202 57
rect 206 49 210 57
rect 214 53 218 57
rect 222 49 226 57
rect 235 49 239 57
rect 248 49 252 57
rect 256 49 260 57
rect 264 49 268 57
rect 272 53 276 57
rect 280 49 284 57
rect 293 49 297 57
rect 301 49 305 57
rect 309 49 313 57
rect 317 49 321 57
rect 330 49 334 57
rect 338 49 342 57
rect 346 53 350 57
rect 354 49 358 57
rect 367 49 371 57
rect 380 49 384 57
rect 388 49 392 57
rect 396 49 400 57
rect 404 53 408 57
rect 412 49 416 57
rect 425 49 429 57
rect 433 49 437 57
rect 441 49 445 57
rect 449 49 453 57
rect 462 49 466 57
rect 470 49 474 57
rect 478 53 482 57
rect 486 49 490 57
rect 499 49 503 57
rect 512 49 516 57
rect 520 49 524 57
rect 528 49 532 57
rect 536 53 540 57
rect 544 49 548 57
rect 557 49 561 57
rect 565 49 569 57
rect 573 49 577 57
<< psubstratepcontact >>
rect 687 911 691 915
rect 715 911 719 915
rect 745 911 749 915
rect 819 911 823 915
rect 847 911 851 915
rect 877 911 881 915
rect 951 911 955 915
rect 979 911 983 915
rect 1009 911 1013 915
rect 1083 911 1087 915
rect 1111 911 1115 915
rect 1141 911 1145 915
rect 347 878 351 882
rect 375 878 379 882
rect 405 878 409 882
rect 668 825 672 829
rect 703 825 707 829
rect 829 825 833 829
rect 853 825 857 829
rect 907 825 914 829
rect 934 825 938 829
rect 988 825 992 829
rect 344 776 348 780
rect 374 776 378 780
rect 402 776 406 780
rect 668 693 672 697
rect 703 693 707 697
rect 829 693 833 697
rect 853 693 857 697
rect 907 693 911 697
rect 934 693 938 697
rect 958 693 962 697
rect 668 561 672 565
rect 703 561 707 565
rect 829 561 833 565
rect 853 561 857 565
rect 907 561 914 565
rect 934 561 938 565
rect 988 561 992 565
rect 1024 561 1028 565
rect 1078 561 1082 565
rect 668 429 672 433
rect 703 429 707 433
rect 829 429 833 433
rect 853 429 857 433
rect 964 429 968 433
rect 215 376 219 380
rect 243 376 247 380
rect 273 376 277 380
rect 347 376 351 380
rect 375 376 379 380
rect 405 376 409 380
rect 479 376 483 380
rect 507 376 511 380
rect 537 376 541 380
rect 986 266 990 270
rect 1014 266 1018 270
rect 1044 266 1048 270
rect 215 236 219 240
rect 243 236 247 240
rect 273 236 277 240
rect 347 236 351 240
rect 375 236 379 240
rect 405 236 409 240
rect 479 236 483 240
rect 507 236 511 240
rect 537 236 541 240
rect 986 180 990 184
rect 1014 180 1018 184
rect 1044 180 1048 184
rect 215 150 219 154
rect 243 150 247 154
rect 273 150 277 154
rect 347 150 351 154
rect 375 150 379 154
rect 405 150 409 154
rect 479 150 483 154
rect 507 150 511 154
rect 537 150 541 154
rect 215 10 219 14
rect 243 10 247 14
rect 273 10 277 14
rect 347 10 351 14
rect 375 10 379 14
rect 405 10 409 14
rect 479 10 483 14
rect 507 10 511 14
rect 537 10 541 14
<< nsubstratencontact >>
rect 687 968 691 972
rect 715 968 719 972
rect 745 968 749 972
rect 782 968 786 972
rect 819 968 823 972
rect 847 968 851 972
rect 877 968 881 972
rect 914 968 918 972
rect 951 968 955 972
rect 979 968 983 972
rect 1009 968 1013 972
rect 1046 968 1050 972
rect 1083 968 1087 972
rect 1111 968 1115 972
rect 1141 968 1145 972
rect 1178 968 1182 972
rect 347 935 351 939
rect 375 935 379 939
rect 405 935 409 939
rect 442 935 446 939
rect 677 891 681 895
rect 706 891 710 895
rect 731 891 735 895
rect 773 891 777 895
rect 829 891 833 895
rect 853 891 857 895
rect 907 891 911 895
rect 934 891 938 895
rect 988 891 992 895
rect 307 833 311 837
rect 344 833 348 837
rect 374 833 378 837
rect 402 833 406 837
rect 677 759 681 763
rect 706 759 710 763
rect 731 759 735 763
rect 773 759 777 763
rect 829 759 833 763
rect 853 759 857 763
rect 907 759 911 763
rect 934 759 938 763
rect 996 759 1000 763
rect 677 627 681 631
rect 706 627 710 631
rect 731 627 735 631
rect 773 627 777 631
rect 829 627 833 631
rect 853 627 857 631
rect 907 627 911 631
rect 934 627 938 631
rect 988 627 992 631
rect 996 627 1000 631
rect 1024 627 1028 631
rect 1078 627 1082 631
rect 677 495 681 499
rect 706 495 710 499
rect 731 495 735 499
rect 773 495 777 499
rect 829 495 833 499
rect 853 495 857 499
rect 907 495 911 499
rect 934 495 938 499
rect 1024 495 1028 499
rect 215 433 219 437
rect 243 433 247 437
rect 273 433 277 437
rect 310 433 314 437
rect 347 433 351 437
rect 375 433 379 437
rect 405 433 409 437
rect 442 433 446 437
rect 479 433 483 437
rect 507 433 511 437
rect 537 433 541 437
rect 574 433 578 437
rect 677 363 681 367
rect 706 363 710 367
rect 731 363 735 367
rect 773 363 777 367
rect 853 363 857 367
rect 907 363 911 367
rect 938 363 942 367
rect 967 363 971 367
rect 992 363 996 367
rect 1034 363 1038 367
rect 986 323 990 327
rect 1014 323 1018 327
rect 1044 323 1048 327
rect 1081 323 1085 327
rect 215 293 219 297
rect 243 293 247 297
rect 273 293 277 297
rect 310 293 314 297
rect 347 293 351 297
rect 375 293 379 297
rect 405 293 409 297
rect 442 293 446 297
rect 479 293 483 297
rect 507 293 511 297
rect 537 293 541 297
rect 574 293 578 297
rect 986 237 990 241
rect 1014 237 1018 241
rect 1044 237 1048 241
rect 1081 237 1085 241
rect 215 207 219 211
rect 243 207 247 211
rect 273 207 277 211
rect 310 207 314 211
rect 347 207 351 211
rect 375 207 379 211
rect 405 207 409 211
rect 442 207 446 211
rect 479 207 483 211
rect 507 207 511 211
rect 537 207 541 211
rect 574 207 578 211
rect 215 67 219 71
rect 243 67 247 71
rect 273 67 277 71
rect 310 67 314 71
rect 347 67 351 71
rect 375 67 379 71
rect 405 67 409 71
rect 442 67 446 71
rect 479 67 483 71
rect 507 67 511 71
rect 537 67 541 71
rect 574 67 578 71
<< polysilicon >>
rect 662 958 664 960
rect 667 958 669 961
rect 683 958 685 960
rect 699 958 701 960
rect 704 958 706 961
rect 725 958 727 961
rect 741 958 743 961
rect 757 958 759 960
rect 762 958 764 961
rect 778 958 780 960
rect 794 958 796 960
rect 799 958 801 961
rect 815 958 817 960
rect 831 958 833 960
rect 836 958 838 961
rect 857 958 859 961
rect 873 958 875 961
rect 889 958 891 960
rect 894 958 896 961
rect 910 958 912 960
rect 926 958 928 960
rect 931 958 933 961
rect 947 958 949 960
rect 963 958 965 960
rect 968 958 970 961
rect 989 958 991 961
rect 1005 958 1007 961
rect 1021 958 1023 960
rect 1026 958 1028 961
rect 1042 958 1044 960
rect 1058 958 1060 960
rect 1063 958 1065 961
rect 1079 958 1081 960
rect 1095 958 1097 960
rect 1100 958 1102 961
rect 1121 958 1123 961
rect 1137 958 1139 961
rect 1153 958 1155 960
rect 1158 958 1160 961
rect 1174 958 1176 960
rect 662 945 664 950
rect 667 948 669 950
rect 662 931 664 941
rect 667 931 669 938
rect 683 931 685 950
rect 699 941 701 950
rect 704 948 706 950
rect 725 948 727 950
rect 741 947 743 950
rect 699 931 701 934
rect 704 931 706 933
rect 725 931 727 933
rect 741 931 743 943
rect 757 941 759 950
rect 762 948 764 950
rect 778 942 780 950
rect 794 945 796 950
rect 799 948 801 950
rect 757 931 759 934
rect 762 931 764 933
rect 778 931 780 938
rect 794 931 796 941
rect 799 931 801 938
rect 815 931 817 950
rect 831 941 833 950
rect 836 948 838 950
rect 857 948 859 950
rect 873 947 875 950
rect 831 931 833 934
rect 836 931 838 933
rect 857 931 859 933
rect 873 931 875 943
rect 889 941 891 950
rect 894 948 896 950
rect 910 942 912 950
rect 926 945 928 950
rect 931 948 933 950
rect 889 931 891 934
rect 894 931 896 933
rect 910 931 912 938
rect 926 931 928 941
rect 931 931 933 938
rect 947 931 949 950
rect 963 941 965 950
rect 968 948 970 950
rect 989 948 991 950
rect 1005 947 1007 950
rect 963 931 965 934
rect 968 931 970 933
rect 989 931 991 933
rect 1005 931 1007 943
rect 1021 941 1023 950
rect 1026 948 1028 950
rect 1042 942 1044 950
rect 1058 945 1060 950
rect 1063 948 1065 950
rect 1021 931 1023 934
rect 1026 931 1028 933
rect 1042 931 1044 938
rect 1058 931 1060 941
rect 1063 931 1065 938
rect 1079 931 1081 950
rect 1095 941 1097 950
rect 1100 948 1102 950
rect 1121 948 1123 950
rect 1137 947 1139 950
rect 1095 931 1097 934
rect 1100 931 1102 933
rect 1121 931 1123 933
rect 1137 931 1139 943
rect 1153 941 1155 950
rect 1158 948 1160 950
rect 1174 942 1176 950
rect 1153 931 1155 934
rect 1158 931 1160 933
rect 1174 931 1176 938
rect 322 925 324 927
rect 327 925 329 928
rect 343 925 345 927
rect 359 925 361 927
rect 364 925 366 928
rect 385 925 387 928
rect 401 925 403 928
rect 417 925 419 927
rect 422 925 424 928
rect 438 925 440 927
rect 662 925 664 927
rect 667 924 669 927
rect 683 925 685 927
rect 699 925 701 927
rect 704 922 706 927
rect 725 922 727 927
rect 741 925 743 927
rect 757 925 759 927
rect 762 922 764 927
rect 778 925 780 927
rect 794 925 796 927
rect 799 924 801 927
rect 815 925 817 927
rect 831 925 833 927
rect 836 922 838 927
rect 857 922 859 927
rect 873 925 875 927
rect 889 925 891 927
rect 894 922 896 927
rect 910 925 912 927
rect 926 925 928 927
rect 931 924 933 927
rect 947 925 949 927
rect 963 925 965 927
rect 968 922 970 927
rect 989 922 991 927
rect 1005 925 1007 927
rect 1021 925 1023 927
rect 1026 922 1028 927
rect 1042 925 1044 927
rect 1058 925 1060 927
rect 1063 924 1065 927
rect 1079 925 1081 927
rect 1095 925 1097 927
rect 1100 922 1102 927
rect 1121 922 1123 927
rect 1137 925 1139 927
rect 1153 925 1155 927
rect 1158 922 1160 927
rect 1174 925 1176 927
rect 322 912 324 917
rect 327 915 329 917
rect 322 898 324 908
rect 327 898 329 905
rect 343 898 345 917
rect 359 908 361 917
rect 364 915 366 917
rect 385 915 387 917
rect 401 914 403 917
rect 359 898 361 901
rect 364 898 366 900
rect 385 898 387 900
rect 401 898 403 910
rect 417 908 419 917
rect 422 915 424 917
rect 417 898 419 901
rect 422 898 424 900
rect 438 898 440 917
rect 322 892 324 894
rect 327 891 329 894
rect 343 892 345 894
rect 359 892 361 894
rect 364 889 366 894
rect 385 889 387 894
rect 401 892 403 894
rect 417 892 419 894
rect 422 889 424 894
rect 438 892 440 894
rect 841 887 843 889
rect 683 881 685 884
rect 727 881 729 884
rect 753 881 755 884
rect 799 881 801 884
rect 753 877 754 881
rect 867 881 869 885
rect 895 887 897 889
rect 922 887 924 889
rect 872 881 874 884
rect 667 874 669 876
rect 683 874 685 877
rect 699 874 701 876
rect 722 874 724 876
rect 727 874 729 877
rect 753 874 755 877
rect 774 874 776 877
rect 794 874 796 876
rect 799 874 801 877
rect 817 874 819 876
rect 446 861 448 864
rect 446 855 448 857
rect 329 852 331 855
rect 667 852 669 866
rect 683 864 685 866
rect 683 852 685 854
rect 699 852 701 866
rect 722 861 724 866
rect 727 864 729 866
rect 753 864 755 866
rect 718 857 724 861
rect 722 852 724 857
rect 727 852 729 854
rect 753 852 755 854
rect 774 852 776 866
rect 794 861 796 866
rect 799 864 801 866
rect 790 857 796 861
rect 794 852 796 857
rect 799 852 801 854
rect 817 852 819 866
rect 841 865 843 879
rect 948 881 950 885
rect 976 887 978 889
rect 953 881 955 884
rect 867 870 869 873
rect 872 871 874 873
rect 868 866 869 870
rect 867 861 869 866
rect 872 861 874 863
rect 841 859 843 861
rect 895 857 897 879
rect 922 865 924 879
rect 948 870 950 873
rect 953 871 955 873
rect 949 866 950 870
rect 948 861 950 866
rect 953 861 955 863
rect 922 859 924 861
rect 976 857 978 879
rect 867 855 869 857
rect 872 852 874 857
rect 948 855 950 857
rect 895 851 897 853
rect 953 852 955 857
rect 976 851 978 853
rect 329 846 331 848
rect 667 846 669 848
rect 683 844 685 848
rect 699 846 701 848
rect 722 846 724 848
rect 684 840 685 844
rect 727 843 729 848
rect 753 844 755 848
rect 774 846 776 848
rect 794 846 796 848
rect 683 837 685 840
rect 728 839 729 843
rect 754 840 755 844
rect 799 843 801 848
rect 817 846 819 848
rect 727 837 729 839
rect 753 836 755 840
rect 800 839 801 843
rect 799 837 801 839
rect 313 823 315 825
rect 329 823 331 826
rect 334 823 336 825
rect 350 823 352 826
rect 366 823 368 826
rect 387 823 389 826
rect 392 823 394 825
rect 408 823 410 825
rect 424 823 426 826
rect 429 823 431 825
rect 313 796 315 815
rect 329 813 331 815
rect 334 806 336 815
rect 350 812 352 815
rect 366 813 368 815
rect 387 813 389 815
rect 329 796 331 798
rect 334 796 336 799
rect 350 796 352 808
rect 392 806 394 815
rect 366 796 368 798
rect 387 796 389 798
rect 392 796 394 799
rect 408 796 410 815
rect 424 813 426 815
rect 429 810 431 815
rect 683 814 685 817
rect 727 815 729 817
rect 684 810 685 814
rect 728 811 729 815
rect 753 814 755 818
rect 799 815 801 817
rect 667 806 669 808
rect 683 806 685 810
rect 699 806 701 808
rect 722 806 724 808
rect 727 806 729 811
rect 754 810 755 814
rect 800 811 801 815
rect 753 806 755 810
rect 774 806 776 808
rect 794 806 796 808
rect 799 806 801 811
rect 817 806 819 808
rect 424 796 426 803
rect 429 796 431 806
rect 867 805 869 808
rect 872 805 874 808
rect 948 805 950 808
rect 953 805 955 808
rect 313 790 315 792
rect 329 787 331 792
rect 334 790 336 792
rect 350 790 352 792
rect 366 787 368 792
rect 387 787 389 792
rect 392 790 394 792
rect 408 790 410 792
rect 424 789 426 792
rect 429 790 431 792
rect 667 788 669 802
rect 683 800 685 802
rect 683 788 685 790
rect 699 788 701 802
rect 722 797 724 802
rect 727 800 729 802
rect 753 800 755 802
rect 718 793 724 797
rect 722 788 724 793
rect 727 788 729 790
rect 753 788 755 790
rect 774 788 776 802
rect 794 797 796 802
rect 799 800 801 802
rect 790 793 796 797
rect 794 788 796 793
rect 799 788 801 790
rect 817 788 819 802
rect 867 789 869 801
rect 872 799 874 801
rect 872 789 874 791
rect 948 789 950 801
rect 953 799 955 801
rect 953 789 955 791
rect 667 778 669 780
rect 683 777 685 780
rect 699 778 701 780
rect 722 778 724 780
rect 727 777 729 780
rect 753 777 755 780
rect 774 777 776 780
rect 794 778 796 780
rect 799 777 801 780
rect 817 778 819 780
rect 867 779 869 781
rect 753 773 754 777
rect 872 776 874 781
rect 948 779 950 781
rect 953 776 955 781
rect 683 770 685 773
rect 727 770 729 773
rect 753 770 755 773
rect 799 770 801 773
rect 683 749 685 752
rect 727 749 729 752
rect 753 749 755 752
rect 799 749 801 752
rect 867 749 869 753
rect 895 755 897 757
rect 946 755 948 757
rect 872 749 874 752
rect 753 745 754 749
rect 667 742 669 744
rect 683 742 685 745
rect 699 742 701 744
rect 722 742 724 744
rect 727 742 729 745
rect 753 742 755 745
rect 774 742 776 745
rect 794 742 796 744
rect 799 742 801 745
rect 817 742 819 744
rect 972 749 974 753
rect 1000 755 1002 757
rect 977 749 979 752
rect 867 738 869 741
rect 872 739 874 741
rect 868 734 869 738
rect 667 720 669 734
rect 683 732 685 734
rect 683 720 685 722
rect 699 720 701 734
rect 722 729 724 734
rect 727 732 729 734
rect 753 732 755 734
rect 718 725 724 729
rect 722 720 724 725
rect 727 720 729 722
rect 753 720 755 722
rect 774 720 776 734
rect 794 729 796 734
rect 799 732 801 734
rect 790 725 796 729
rect 794 720 796 725
rect 799 720 801 722
rect 817 720 819 734
rect 867 729 869 734
rect 872 729 874 731
rect 895 725 897 747
rect 946 733 948 747
rect 972 738 974 741
rect 977 739 979 741
rect 973 734 974 738
rect 972 729 974 734
rect 977 729 979 731
rect 946 727 948 729
rect 1000 725 1002 747
rect 867 723 869 725
rect 872 720 874 725
rect 972 723 974 725
rect 895 719 897 721
rect 977 720 979 725
rect 1000 719 1002 721
rect 667 714 669 716
rect 683 712 685 716
rect 699 714 701 716
rect 722 714 724 716
rect 684 708 685 712
rect 727 711 729 716
rect 753 712 755 716
rect 774 714 776 716
rect 794 714 796 716
rect 683 705 685 708
rect 728 707 729 711
rect 754 708 755 712
rect 799 711 801 716
rect 817 714 819 716
rect 727 705 729 707
rect 753 704 755 708
rect 800 707 801 711
rect 799 705 801 707
rect 683 682 685 685
rect 727 683 729 685
rect 684 678 685 682
rect 728 679 729 683
rect 753 682 755 686
rect 799 683 801 685
rect 667 674 669 676
rect 683 674 685 678
rect 699 674 701 676
rect 722 674 724 676
rect 727 674 729 679
rect 754 678 755 682
rect 800 679 801 683
rect 753 674 755 678
rect 774 674 776 676
rect 794 674 796 676
rect 799 674 801 679
rect 817 674 819 676
rect 867 674 869 677
rect 872 674 874 677
rect 972 674 974 677
rect 977 674 979 677
rect 667 656 669 670
rect 683 668 685 670
rect 683 656 685 658
rect 699 656 701 670
rect 722 665 724 670
rect 727 668 729 670
rect 753 668 755 670
rect 718 661 724 665
rect 722 656 724 661
rect 727 656 729 658
rect 753 656 755 658
rect 774 656 776 670
rect 794 665 796 670
rect 799 668 801 670
rect 790 661 796 665
rect 794 656 796 661
rect 799 656 801 658
rect 817 656 819 670
rect 867 658 869 670
rect 872 668 874 670
rect 872 658 874 660
rect 972 658 974 670
rect 977 668 979 670
rect 977 658 979 660
rect 867 648 869 650
rect 667 646 669 648
rect 683 645 685 648
rect 699 646 701 648
rect 722 646 724 648
rect 727 645 729 648
rect 753 645 755 648
rect 774 645 776 648
rect 794 646 796 648
rect 799 645 801 648
rect 817 646 819 648
rect 872 645 874 650
rect 972 648 974 650
rect 977 645 979 650
rect 753 641 754 645
rect 683 638 685 641
rect 727 638 729 641
rect 753 638 755 641
rect 799 638 801 641
rect 683 617 685 620
rect 727 617 729 620
rect 753 617 755 620
rect 799 617 801 620
rect 867 617 869 621
rect 895 623 897 625
rect 922 623 924 625
rect 872 617 874 620
rect 753 613 754 617
rect 667 610 669 612
rect 683 610 685 613
rect 699 610 701 612
rect 722 610 724 612
rect 727 610 729 613
rect 753 610 755 613
rect 774 610 776 613
rect 794 610 796 612
rect 799 610 801 613
rect 817 610 819 612
rect 948 617 950 621
rect 976 623 978 625
rect 1012 623 1014 625
rect 953 617 955 620
rect 867 606 869 609
rect 872 607 874 609
rect 868 602 869 606
rect 667 588 669 602
rect 683 600 685 602
rect 683 588 685 590
rect 699 588 701 602
rect 722 597 724 602
rect 727 600 729 602
rect 753 600 755 602
rect 718 593 724 597
rect 722 588 724 593
rect 727 588 729 590
rect 753 588 755 590
rect 774 588 776 602
rect 794 597 796 602
rect 799 600 801 602
rect 790 593 796 597
rect 794 588 796 593
rect 799 588 801 590
rect 817 588 819 602
rect 867 597 869 602
rect 872 597 874 599
rect 895 593 897 615
rect 922 601 924 615
rect 1038 617 1040 621
rect 1066 623 1068 625
rect 1043 617 1045 620
rect 948 606 950 609
rect 953 607 955 609
rect 949 602 950 606
rect 948 597 950 602
rect 953 597 955 599
rect 922 595 924 597
rect 976 593 978 615
rect 1012 601 1014 615
rect 1038 606 1040 609
rect 1043 607 1045 609
rect 1039 602 1040 606
rect 1038 597 1040 602
rect 1043 597 1045 599
rect 1012 595 1014 597
rect 1066 593 1068 615
rect 867 591 869 593
rect 872 588 874 593
rect 948 591 950 593
rect 895 587 897 589
rect 953 588 955 593
rect 1038 591 1040 593
rect 976 587 978 589
rect 1043 588 1045 593
rect 1066 587 1068 589
rect 667 582 669 584
rect 683 580 685 584
rect 699 582 701 584
rect 722 582 724 584
rect 684 576 685 580
rect 727 579 729 584
rect 753 580 755 584
rect 774 582 776 584
rect 794 582 796 584
rect 683 573 685 576
rect 728 575 729 579
rect 754 576 755 580
rect 799 579 801 584
rect 817 582 819 584
rect 727 573 729 575
rect 753 572 755 576
rect 800 575 801 579
rect 799 573 801 575
rect 683 550 685 553
rect 727 551 729 553
rect 684 546 685 550
rect 728 547 729 551
rect 753 550 755 554
rect 799 551 801 553
rect 667 542 669 544
rect 683 542 685 546
rect 699 542 701 544
rect 722 542 724 544
rect 727 542 729 547
rect 754 546 755 550
rect 800 547 801 551
rect 753 542 755 546
rect 774 542 776 544
rect 794 542 796 544
rect 799 542 801 547
rect 817 542 819 544
rect 867 539 869 542
rect 872 539 874 542
rect 948 539 950 542
rect 953 539 955 542
rect 1038 539 1040 542
rect 1043 539 1045 542
rect 667 524 669 538
rect 683 536 685 538
rect 683 524 685 526
rect 699 524 701 538
rect 722 533 724 538
rect 727 536 729 538
rect 753 536 755 538
rect 718 529 724 533
rect 722 524 724 529
rect 727 524 729 526
rect 753 524 755 526
rect 774 524 776 538
rect 794 533 796 538
rect 799 536 801 538
rect 790 529 796 533
rect 794 524 796 529
rect 799 524 801 526
rect 817 524 819 538
rect 867 523 869 535
rect 872 533 874 535
rect 872 523 874 525
rect 948 523 950 535
rect 953 533 955 535
rect 953 523 955 525
rect 1038 523 1040 535
rect 1043 533 1045 535
rect 1043 523 1045 525
rect 667 514 669 516
rect 683 513 685 516
rect 699 514 701 516
rect 722 514 724 516
rect 727 513 729 516
rect 753 513 755 516
rect 774 513 776 516
rect 794 514 796 516
rect 799 513 801 516
rect 817 514 819 516
rect 867 513 869 515
rect 753 509 754 513
rect 872 510 874 515
rect 948 513 950 515
rect 953 510 955 515
rect 1038 513 1040 515
rect 1043 510 1045 515
rect 683 506 685 509
rect 727 506 729 509
rect 753 506 755 509
rect 799 506 801 509
rect 683 485 685 488
rect 727 485 729 488
rect 753 485 755 488
rect 799 485 801 488
rect 867 485 869 489
rect 895 491 897 493
rect 872 485 874 488
rect 753 481 754 485
rect 667 478 669 480
rect 683 478 685 481
rect 699 478 701 480
rect 722 478 724 480
rect 727 478 729 481
rect 753 478 755 481
rect 774 478 776 481
rect 794 478 796 480
rect 799 478 801 481
rect 817 478 819 480
rect 867 474 869 477
rect 872 475 874 477
rect 868 470 869 474
rect 667 456 669 470
rect 683 468 685 470
rect 683 456 685 458
rect 699 456 701 470
rect 722 465 724 470
rect 727 468 729 470
rect 753 468 755 470
rect 718 461 724 465
rect 722 456 724 461
rect 727 456 729 458
rect 753 456 755 458
rect 774 456 776 470
rect 794 465 796 470
rect 799 468 801 470
rect 790 461 796 465
rect 794 456 796 461
rect 799 456 801 458
rect 817 456 819 470
rect 867 465 869 470
rect 872 465 874 467
rect 895 461 897 483
rect 867 459 869 461
rect 872 456 874 461
rect 895 455 897 457
rect 667 450 669 452
rect 683 448 685 452
rect 699 450 701 452
rect 722 450 724 452
rect 684 444 685 448
rect 727 447 729 452
rect 753 448 755 452
rect 774 450 776 452
rect 794 450 796 452
rect 683 441 685 444
rect 728 443 729 447
rect 754 444 755 448
rect 799 447 801 452
rect 817 450 819 452
rect 727 441 729 443
rect 753 440 755 444
rect 800 443 801 447
rect 799 441 801 443
rect 190 423 192 425
rect 195 423 197 426
rect 211 423 213 425
rect 227 423 229 425
rect 232 423 234 426
rect 253 423 255 426
rect 269 423 271 426
rect 285 423 287 425
rect 290 423 292 426
rect 306 423 308 425
rect 322 423 324 425
rect 327 423 329 426
rect 343 423 345 425
rect 359 423 361 425
rect 364 423 366 426
rect 385 423 387 426
rect 401 423 403 426
rect 417 423 419 425
rect 422 423 424 426
rect 438 423 440 425
rect 454 423 456 425
rect 459 423 461 426
rect 475 423 477 425
rect 491 423 493 425
rect 496 423 498 426
rect 517 423 519 426
rect 533 423 535 426
rect 549 423 551 425
rect 554 423 556 426
rect 570 423 572 425
rect 683 418 685 421
rect 727 419 729 421
rect 190 410 192 415
rect 195 413 197 415
rect 190 396 192 406
rect 195 396 197 403
rect 211 396 213 415
rect 227 406 229 415
rect 232 413 234 415
rect 253 413 255 415
rect 269 412 271 415
rect 227 396 229 399
rect 232 396 234 398
rect 253 396 255 398
rect 269 396 271 408
rect 285 406 287 415
rect 290 413 292 415
rect 285 396 287 399
rect 290 396 292 398
rect 306 396 308 415
rect 322 412 324 415
rect 327 413 329 415
rect 322 396 324 408
rect 327 396 329 403
rect 343 396 345 415
rect 359 406 361 415
rect 364 413 366 415
rect 385 413 387 415
rect 401 412 403 415
rect 359 396 361 399
rect 364 396 366 398
rect 385 396 387 398
rect 401 396 403 408
rect 417 406 419 415
rect 422 413 424 415
rect 417 396 419 399
rect 422 396 424 398
rect 438 396 440 415
rect 454 412 456 415
rect 459 413 461 415
rect 454 396 456 408
rect 459 396 461 403
rect 475 396 477 415
rect 491 406 493 415
rect 496 413 498 415
rect 517 413 519 415
rect 533 412 535 415
rect 491 396 493 399
rect 496 396 498 398
rect 517 396 519 398
rect 533 396 535 408
rect 549 406 551 415
rect 554 413 556 415
rect 570 407 572 415
rect 684 414 685 418
rect 728 415 729 419
rect 753 418 755 422
rect 799 419 801 421
rect 667 410 669 412
rect 683 410 685 414
rect 699 410 701 412
rect 722 410 724 412
rect 727 410 729 415
rect 754 414 755 418
rect 800 415 801 419
rect 944 418 946 421
rect 988 419 990 421
rect 753 410 755 414
rect 774 410 776 412
rect 794 410 796 412
rect 799 410 801 415
rect 945 414 946 418
rect 989 415 990 419
rect 1014 418 1016 422
rect 1060 419 1062 421
rect 817 410 819 412
rect 901 410 903 413
rect 919 410 921 413
rect 944 410 946 414
rect 960 410 962 412
rect 983 410 985 412
rect 988 410 990 415
rect 1015 414 1016 418
rect 1061 415 1062 419
rect 1014 410 1016 414
rect 1035 410 1037 412
rect 1055 410 1057 412
rect 1060 410 1062 415
rect 1078 410 1080 412
rect 549 396 551 399
rect 554 396 556 398
rect 570 396 572 403
rect 667 392 669 406
rect 683 404 685 406
rect 683 392 685 394
rect 699 392 701 406
rect 722 401 724 406
rect 727 404 729 406
rect 753 404 755 406
rect 718 397 724 401
rect 722 392 724 397
rect 727 392 729 394
rect 753 392 755 394
rect 774 392 776 406
rect 794 401 796 406
rect 799 404 801 406
rect 790 397 796 401
rect 794 392 796 397
rect 799 392 801 394
rect 817 392 819 406
rect 867 403 869 406
rect 872 403 874 406
rect 901 401 903 406
rect 190 390 192 392
rect 195 389 197 392
rect 211 390 213 392
rect 227 390 229 392
rect 232 387 234 392
rect 253 387 255 392
rect 269 390 271 392
rect 285 390 287 392
rect 290 387 292 392
rect 306 390 308 392
rect 322 390 324 392
rect 327 389 329 392
rect 343 390 345 392
rect 359 390 361 392
rect 364 387 366 392
rect 385 387 387 392
rect 401 390 403 392
rect 417 390 419 392
rect 422 387 424 392
rect 438 390 440 392
rect 454 390 456 392
rect 459 389 461 392
rect 475 390 477 392
rect 491 390 493 392
rect 496 387 498 392
rect 517 387 519 392
rect 533 390 535 392
rect 549 390 551 392
rect 554 387 556 392
rect 570 390 572 392
rect 867 387 869 399
rect 872 397 874 399
rect 901 392 903 397
rect 919 392 921 406
rect 944 404 946 406
rect 944 392 946 394
rect 960 392 962 406
rect 983 401 985 406
rect 988 404 990 406
rect 1014 404 1016 406
rect 979 397 985 401
rect 983 392 985 397
rect 988 392 990 394
rect 1014 392 1016 394
rect 1035 392 1037 406
rect 1055 401 1057 406
rect 1060 404 1062 406
rect 1051 397 1057 401
rect 1055 392 1057 397
rect 1060 392 1062 394
rect 1078 392 1080 406
rect 872 387 874 389
rect 667 382 669 384
rect 683 381 685 384
rect 699 382 701 384
rect 722 382 724 384
rect 727 381 729 384
rect 753 381 755 384
rect 774 381 776 384
rect 794 382 796 384
rect 799 381 801 384
rect 817 382 819 384
rect 753 377 754 381
rect 901 381 903 384
rect 919 381 921 384
rect 944 381 946 384
rect 960 382 962 384
rect 983 382 985 384
rect 988 381 990 384
rect 1014 381 1016 384
rect 1035 381 1037 384
rect 1055 382 1057 384
rect 1060 381 1062 384
rect 1078 382 1080 384
rect 867 377 869 379
rect 683 374 685 377
rect 727 374 729 377
rect 753 374 755 377
rect 799 374 801 377
rect 872 374 874 379
rect 1014 377 1015 381
rect 944 374 946 377
rect 988 374 990 377
rect 1014 374 1016 377
rect 1060 374 1062 377
rect 305 352 307 355
rect 329 352 331 355
rect 1087 350 1090 352
rect 1094 350 1097 352
rect 305 346 307 348
rect 329 346 331 348
rect 325 341 327 343
rect 325 334 327 337
rect 314 323 316 325
rect 320 323 339 325
rect 305 318 307 320
rect 329 318 331 320
rect 305 311 307 314
rect 329 311 331 314
rect 961 313 963 315
rect 966 313 968 316
rect 982 313 984 315
rect 998 313 1000 315
rect 1003 313 1005 316
rect 1024 313 1026 316
rect 1040 313 1042 316
rect 1056 313 1058 315
rect 1061 313 1063 316
rect 1077 313 1079 315
rect 961 300 963 305
rect 966 303 968 305
rect 961 286 963 296
rect 966 286 968 293
rect 982 286 984 305
rect 998 296 1000 305
rect 1003 303 1005 305
rect 1024 303 1026 305
rect 1040 302 1042 305
rect 998 286 1000 289
rect 1003 286 1005 288
rect 1024 286 1026 288
rect 1040 286 1042 298
rect 1056 296 1058 305
rect 1061 303 1063 305
rect 1056 286 1058 289
rect 1061 286 1063 288
rect 1077 286 1079 305
rect 190 283 192 285
rect 195 283 197 286
rect 211 283 213 285
rect 227 283 229 285
rect 232 283 234 286
rect 253 283 255 286
rect 269 283 271 286
rect 285 283 287 285
rect 290 283 292 286
rect 306 283 308 285
rect 322 283 324 285
rect 327 283 329 286
rect 343 283 345 285
rect 359 283 361 285
rect 364 283 366 286
rect 385 283 387 286
rect 401 283 403 286
rect 417 283 419 285
rect 422 283 424 286
rect 438 283 440 285
rect 454 283 456 285
rect 459 283 461 286
rect 475 283 477 285
rect 491 283 493 285
rect 496 283 498 286
rect 517 283 519 286
rect 533 283 535 286
rect 549 283 551 285
rect 554 283 556 286
rect 570 283 572 285
rect 961 280 963 282
rect 966 279 968 282
rect 982 280 984 282
rect 998 280 1000 282
rect 1003 277 1005 282
rect 1024 277 1026 282
rect 1040 280 1042 282
rect 1056 280 1058 282
rect 1061 277 1063 282
rect 1077 280 1079 282
rect 190 270 192 275
rect 195 273 197 275
rect 190 256 192 266
rect 195 256 197 263
rect 211 256 213 275
rect 227 266 229 275
rect 232 273 234 275
rect 253 273 255 275
rect 269 272 271 275
rect 227 256 229 259
rect 232 256 234 258
rect 253 256 255 258
rect 269 256 271 268
rect 285 266 287 275
rect 290 273 292 275
rect 285 256 287 259
rect 290 256 292 258
rect 306 256 308 275
rect 322 272 324 275
rect 327 273 329 275
rect 322 256 324 268
rect 327 256 329 263
rect 343 256 345 275
rect 359 266 361 275
rect 364 273 366 275
rect 385 273 387 275
rect 401 272 403 275
rect 359 256 361 259
rect 364 256 366 258
rect 385 256 387 258
rect 401 256 403 268
rect 417 266 419 275
rect 422 273 424 275
rect 417 256 419 259
rect 422 256 424 258
rect 438 256 440 275
rect 454 272 456 275
rect 459 273 461 275
rect 454 256 456 268
rect 459 256 461 263
rect 475 256 477 275
rect 491 266 493 275
rect 496 273 498 275
rect 517 273 519 275
rect 533 272 535 275
rect 491 256 493 259
rect 496 256 498 258
rect 517 256 519 258
rect 533 256 535 268
rect 549 266 551 275
rect 554 273 556 275
rect 570 267 572 275
rect 549 256 551 259
rect 554 256 556 258
rect 570 256 572 263
rect 190 250 192 252
rect 195 249 197 252
rect 211 250 213 252
rect 227 250 229 252
rect 232 247 234 252
rect 253 247 255 252
rect 269 250 271 252
rect 285 250 287 252
rect 290 247 292 252
rect 306 250 308 252
rect 322 250 324 252
rect 327 249 329 252
rect 343 250 345 252
rect 359 250 361 252
rect 364 247 366 252
rect 385 247 387 252
rect 401 250 403 252
rect 417 250 419 252
rect 422 247 424 252
rect 438 250 440 252
rect 454 250 456 252
rect 459 249 461 252
rect 475 250 477 252
rect 491 250 493 252
rect 496 247 498 252
rect 517 247 519 252
rect 533 250 535 252
rect 549 250 551 252
rect 554 247 556 252
rect 570 250 572 252
rect 961 227 963 229
rect 966 227 968 230
rect 982 227 984 229
rect 998 227 1000 229
rect 1003 227 1005 230
rect 1024 227 1026 230
rect 1040 227 1042 230
rect 1056 227 1058 229
rect 1061 227 1063 230
rect 1077 227 1079 229
rect 961 214 963 219
rect 966 217 968 219
rect 961 200 963 210
rect 966 200 968 207
rect 982 200 984 219
rect 998 210 1000 219
rect 1003 217 1005 219
rect 1024 217 1026 219
rect 1040 216 1042 219
rect 998 200 1000 203
rect 1003 200 1005 202
rect 1024 200 1026 202
rect 1040 200 1042 212
rect 1056 210 1058 219
rect 1061 217 1063 219
rect 1056 200 1058 203
rect 1061 200 1063 202
rect 1077 200 1079 219
rect 1099 206 1102 208
rect 1106 206 1109 208
rect 190 197 192 199
rect 195 197 197 200
rect 211 197 213 199
rect 227 197 229 199
rect 232 197 234 200
rect 253 197 255 200
rect 269 197 271 200
rect 285 197 287 199
rect 290 197 292 200
rect 306 197 308 199
rect 322 197 324 199
rect 327 197 329 200
rect 343 197 345 199
rect 359 197 361 199
rect 364 197 366 200
rect 385 197 387 200
rect 401 197 403 200
rect 417 197 419 199
rect 422 197 424 200
rect 438 197 440 199
rect 454 197 456 199
rect 459 197 461 200
rect 475 197 477 199
rect 491 197 493 199
rect 496 197 498 200
rect 517 197 519 200
rect 533 197 535 200
rect 549 197 551 199
rect 554 197 556 200
rect 570 197 572 199
rect 961 194 963 196
rect 966 193 968 196
rect 982 194 984 196
rect 998 194 1000 196
rect 1003 191 1005 196
rect 1024 191 1026 196
rect 1040 194 1042 196
rect 1056 194 1058 196
rect 1061 191 1063 196
rect 1077 194 1079 196
rect 190 184 192 189
rect 195 187 197 189
rect 190 170 192 180
rect 195 170 197 177
rect 211 170 213 189
rect 227 180 229 189
rect 232 187 234 189
rect 253 187 255 189
rect 269 186 271 189
rect 227 170 229 173
rect 232 170 234 172
rect 253 170 255 172
rect 269 170 271 182
rect 285 180 287 189
rect 290 187 292 189
rect 285 170 287 173
rect 290 170 292 172
rect 306 170 308 189
rect 322 186 324 189
rect 327 187 329 189
rect 322 170 324 182
rect 327 170 329 177
rect 343 170 345 189
rect 359 180 361 189
rect 364 187 366 189
rect 385 187 387 189
rect 401 186 403 189
rect 359 170 361 173
rect 364 170 366 172
rect 385 170 387 172
rect 401 170 403 182
rect 417 180 419 189
rect 422 187 424 189
rect 417 170 419 173
rect 422 170 424 172
rect 438 170 440 189
rect 454 186 456 189
rect 459 187 461 189
rect 454 170 456 182
rect 459 170 461 177
rect 475 170 477 189
rect 491 180 493 189
rect 496 187 498 189
rect 517 187 519 189
rect 533 186 535 189
rect 491 170 493 173
rect 496 170 498 172
rect 517 170 519 172
rect 533 170 535 182
rect 549 180 551 189
rect 554 187 556 189
rect 570 181 572 189
rect 549 170 551 173
rect 554 170 556 172
rect 570 170 572 177
rect 190 164 192 166
rect 195 163 197 166
rect 211 164 213 166
rect 227 164 229 166
rect 232 161 234 166
rect 253 161 255 166
rect 269 164 271 166
rect 285 164 287 166
rect 290 161 292 166
rect 306 164 308 166
rect 322 164 324 166
rect 327 163 329 166
rect 343 164 345 166
rect 359 164 361 166
rect 364 161 366 166
rect 385 161 387 166
rect 401 164 403 166
rect 417 164 419 166
rect 422 161 424 166
rect 438 164 440 166
rect 454 164 456 166
rect 459 163 461 166
rect 475 164 477 166
rect 491 164 493 166
rect 496 161 498 166
rect 517 161 519 166
rect 533 164 535 166
rect 549 164 551 166
rect 554 161 556 166
rect 570 164 572 166
rect 422 126 424 129
rect 446 126 448 129
rect 422 120 424 122
rect 446 120 448 122
rect 442 115 444 117
rect 442 108 444 111
rect 431 97 433 99
rect 437 97 456 99
rect 422 92 424 94
rect 446 92 448 94
rect 422 85 424 88
rect 446 85 448 88
rect 190 57 192 59
rect 195 57 197 60
rect 211 57 213 59
rect 227 57 229 59
rect 232 57 234 60
rect 253 57 255 60
rect 269 57 271 60
rect 285 57 287 59
rect 290 57 292 60
rect 306 57 308 59
rect 322 57 324 59
rect 327 57 329 60
rect 343 57 345 59
rect 359 57 361 59
rect 364 57 366 60
rect 385 57 387 60
rect 401 57 403 60
rect 417 57 419 59
rect 422 57 424 60
rect 438 57 440 59
rect 454 57 456 59
rect 459 57 461 60
rect 475 57 477 59
rect 491 57 493 59
rect 496 57 498 60
rect 517 57 519 60
rect 533 57 535 60
rect 549 57 551 59
rect 554 57 556 60
rect 570 57 572 59
rect 190 44 192 49
rect 195 47 197 49
rect 190 30 192 40
rect 195 30 197 37
rect 211 30 213 49
rect 227 40 229 49
rect 232 47 234 49
rect 253 47 255 49
rect 269 46 271 49
rect 227 30 229 33
rect 232 30 234 32
rect 253 30 255 32
rect 269 30 271 42
rect 285 40 287 49
rect 290 47 292 49
rect 285 30 287 33
rect 290 30 292 32
rect 306 30 308 49
rect 322 46 324 49
rect 327 47 329 49
rect 322 30 324 42
rect 327 30 329 37
rect 343 30 345 49
rect 359 40 361 49
rect 364 47 366 49
rect 385 47 387 49
rect 401 46 403 49
rect 359 30 361 33
rect 364 30 366 32
rect 385 30 387 32
rect 401 30 403 42
rect 417 40 419 49
rect 422 47 424 49
rect 417 30 419 33
rect 422 30 424 32
rect 438 30 440 49
rect 454 46 456 49
rect 459 47 461 49
rect 454 30 456 42
rect 459 30 461 37
rect 475 30 477 49
rect 491 40 493 49
rect 496 47 498 49
rect 517 47 519 49
rect 533 46 535 49
rect 491 30 493 33
rect 496 30 498 32
rect 517 30 519 32
rect 533 30 535 42
rect 549 40 551 49
rect 554 47 556 49
rect 570 41 572 49
rect 549 30 551 33
rect 554 30 556 32
rect 570 30 572 37
rect 190 24 192 26
rect 195 23 197 26
rect 211 24 213 26
rect 227 24 229 26
rect 232 21 234 26
rect 253 21 255 26
rect 269 24 271 26
rect 285 24 287 26
rect 290 21 292 26
rect 306 24 308 26
rect 322 24 324 26
rect 327 23 329 26
rect 343 24 345 26
rect 359 24 361 26
rect 364 21 366 26
rect 385 21 387 26
rect 401 24 403 26
rect 417 24 419 26
rect 422 21 424 26
rect 438 24 440 26
rect 454 24 456 26
rect 459 23 461 26
rect 475 24 477 26
rect 491 24 493 26
rect 496 21 498 26
rect 517 21 519 26
rect 533 24 535 26
rect 549 24 551 26
rect 554 21 556 26
rect 570 24 572 26
<< polycontact >>
rect 667 961 671 965
rect 704 961 708 965
rect 724 961 728 965
rect 762 961 766 965
rect 799 961 803 965
rect 836 961 840 965
rect 856 961 860 965
rect 894 961 898 965
rect 931 961 935 965
rect 968 961 972 965
rect 988 961 992 965
rect 1026 961 1030 965
rect 1063 961 1067 965
rect 1100 961 1104 965
rect 1120 961 1124 965
rect 1158 961 1162 965
rect 661 941 665 945
rect 679 943 683 947
rect 327 928 331 932
rect 364 928 368 932
rect 384 928 388 932
rect 422 928 426 932
rect 739 943 743 947
rect 697 934 701 941
rect 755 934 759 941
rect 776 938 780 942
rect 793 941 797 945
rect 811 943 815 947
rect 871 943 875 947
rect 829 934 833 941
rect 887 934 891 941
rect 908 938 912 942
rect 925 941 929 945
rect 943 943 947 947
rect 1003 943 1007 947
rect 961 934 965 941
rect 1019 934 1023 941
rect 1040 938 1044 942
rect 1057 941 1061 945
rect 1075 943 1079 947
rect 1135 943 1139 947
rect 1093 934 1097 941
rect 1151 934 1155 941
rect 1172 938 1176 942
rect 667 920 671 924
rect 704 918 708 922
rect 724 918 728 922
rect 760 918 764 922
rect 799 920 803 924
rect 836 918 840 922
rect 856 918 860 922
rect 892 918 896 922
rect 931 920 935 924
rect 968 918 972 922
rect 988 918 992 922
rect 1024 918 1028 922
rect 1063 920 1067 924
rect 1100 918 1104 922
rect 1120 918 1124 922
rect 1156 918 1160 922
rect 321 908 325 912
rect 339 910 343 914
rect 399 910 403 914
rect 357 901 361 908
rect 415 901 419 908
rect 434 905 438 909
rect 327 887 331 891
rect 364 885 368 889
rect 384 885 388 889
rect 420 885 424 889
rect 683 877 687 881
rect 727 877 731 881
rect 754 877 758 881
rect 799 877 803 881
rect 872 884 876 888
rect 445 864 449 868
rect 837 870 841 874
rect 328 855 332 859
rect 663 857 667 861
rect 695 858 699 862
rect 714 857 718 861
rect 770 858 774 862
rect 786 857 790 861
rect 813 857 817 861
rect 953 884 957 888
rect 864 866 868 870
rect 891 862 895 866
rect 918 870 922 874
rect 945 866 949 870
rect 972 862 976 866
rect 870 848 874 852
rect 951 848 955 852
rect 680 840 684 844
rect 724 839 728 843
rect 749 840 754 844
rect 796 839 800 843
rect 327 826 331 830
rect 365 826 369 830
rect 385 826 389 830
rect 422 826 426 830
rect 315 803 319 807
rect 350 808 354 812
rect 334 799 338 806
rect 392 799 396 806
rect 410 808 414 812
rect 680 810 684 814
rect 724 811 728 815
rect 428 806 432 810
rect 749 810 754 814
rect 796 811 800 815
rect 872 808 876 812
rect 953 808 957 812
rect 663 793 667 797
rect 329 783 333 787
rect 365 783 369 787
rect 385 783 389 787
rect 422 785 426 789
rect 695 792 699 796
rect 714 793 718 797
rect 770 792 774 796
rect 786 793 790 797
rect 813 793 817 797
rect 861 792 867 796
rect 942 792 948 796
rect 683 773 687 777
rect 727 773 731 777
rect 754 773 758 777
rect 799 773 803 777
rect 870 772 874 776
rect 951 772 955 776
rect 872 752 876 756
rect 683 745 687 749
rect 727 745 731 749
rect 754 745 758 749
rect 799 745 803 749
rect 977 752 981 756
rect 864 734 868 738
rect 663 725 667 729
rect 695 726 699 730
rect 714 725 718 729
rect 770 726 774 730
rect 786 725 790 729
rect 813 725 817 729
rect 891 730 895 734
rect 942 738 946 742
rect 969 734 973 738
rect 996 730 1000 734
rect 870 716 874 720
rect 975 716 979 720
rect 680 708 684 712
rect 724 707 728 711
rect 749 708 754 712
rect 796 707 800 711
rect 680 678 684 682
rect 724 679 728 683
rect 749 678 754 682
rect 796 679 800 683
rect 872 677 876 681
rect 977 677 981 681
rect 663 661 667 665
rect 695 660 699 664
rect 714 661 718 665
rect 770 660 774 664
rect 786 661 790 665
rect 813 661 817 665
rect 861 661 867 665
rect 966 661 972 665
rect 683 641 687 645
rect 727 641 731 645
rect 754 641 758 645
rect 799 641 803 645
rect 870 641 874 645
rect 975 641 979 645
rect 872 620 876 624
rect 683 613 687 617
rect 727 613 731 617
rect 754 613 758 617
rect 799 613 803 617
rect 953 620 957 624
rect 864 602 868 606
rect 663 593 667 597
rect 695 594 699 598
rect 714 593 718 597
rect 770 594 774 598
rect 786 593 790 597
rect 813 593 817 597
rect 891 598 895 602
rect 918 606 922 610
rect 1043 620 1047 624
rect 945 602 949 606
rect 972 598 976 602
rect 1008 606 1012 610
rect 1035 602 1039 606
rect 1062 598 1066 602
rect 870 584 874 588
rect 951 584 955 588
rect 1041 584 1045 588
rect 680 576 684 580
rect 724 575 728 579
rect 749 576 754 580
rect 796 575 800 579
rect 680 546 684 550
rect 724 547 728 551
rect 749 546 754 550
rect 796 547 800 551
rect 872 542 876 546
rect 953 542 957 546
rect 1043 542 1047 546
rect 663 529 667 533
rect 695 528 699 532
rect 714 529 718 533
rect 770 528 774 532
rect 786 529 790 533
rect 813 529 817 533
rect 861 526 867 530
rect 942 526 948 530
rect 1032 526 1038 530
rect 683 509 687 513
rect 727 509 731 513
rect 754 509 758 513
rect 799 509 803 513
rect 870 506 874 510
rect 951 506 955 510
rect 1041 506 1045 510
rect 872 488 876 492
rect 683 481 687 485
rect 727 481 731 485
rect 754 481 758 485
rect 799 481 803 485
rect 864 470 868 474
rect 663 461 667 465
rect 695 462 699 466
rect 714 461 718 465
rect 770 462 774 466
rect 786 461 790 465
rect 813 461 817 465
rect 891 466 895 470
rect 870 452 874 456
rect 680 444 684 448
rect 724 443 728 447
rect 749 444 754 448
rect 796 443 800 447
rect 195 426 199 430
rect 232 426 236 430
rect 252 426 256 430
rect 290 426 294 430
rect 327 426 331 430
rect 364 426 368 430
rect 384 426 388 430
rect 422 426 426 430
rect 459 426 463 430
rect 496 426 500 430
rect 516 426 520 430
rect 554 426 558 430
rect 189 406 193 410
rect 207 408 211 412
rect 267 408 271 412
rect 225 399 229 406
rect 283 399 287 406
rect 302 403 306 407
rect 320 408 324 412
rect 339 408 343 412
rect 399 408 403 412
rect 357 399 361 406
rect 415 399 419 406
rect 434 403 438 407
rect 452 408 456 412
rect 471 408 475 412
rect 531 408 535 412
rect 489 399 493 406
rect 680 414 684 418
rect 724 415 728 419
rect 749 414 754 418
rect 796 415 800 419
rect 941 414 945 418
rect 985 415 989 419
rect 1010 414 1015 418
rect 1057 415 1061 419
rect 547 399 551 406
rect 568 403 572 407
rect 872 406 876 410
rect 663 397 667 401
rect 695 396 699 400
rect 714 397 718 401
rect 770 396 774 400
rect 786 397 790 401
rect 813 397 817 401
rect 195 385 199 389
rect 232 383 236 387
rect 252 383 256 387
rect 288 383 292 387
rect 327 385 331 389
rect 364 383 368 387
rect 384 383 388 387
rect 420 383 424 387
rect 459 385 463 389
rect 496 383 500 387
rect 516 383 520 387
rect 552 383 556 387
rect 861 390 867 394
rect 899 397 903 401
rect 956 396 960 400
rect 975 397 979 401
rect 1031 396 1035 400
rect 1047 397 1051 401
rect 1074 397 1078 401
rect 683 377 687 381
rect 727 377 731 381
rect 754 377 758 381
rect 799 377 803 381
rect 944 377 948 381
rect 988 377 992 381
rect 1015 377 1019 381
rect 1060 377 1064 381
rect 870 370 874 374
rect 304 355 308 359
rect 328 355 332 359
rect 1083 349 1087 353
rect 324 330 328 334
rect 339 322 343 326
rect 966 316 970 320
rect 1003 316 1007 320
rect 1023 316 1027 320
rect 1061 316 1065 320
rect 304 307 308 311
rect 328 307 332 311
rect 960 296 964 300
rect 978 298 982 302
rect 195 286 199 290
rect 232 286 236 290
rect 252 286 256 290
rect 290 286 294 290
rect 327 286 331 290
rect 364 286 368 290
rect 384 286 388 290
rect 422 286 426 290
rect 459 286 463 290
rect 496 286 500 290
rect 516 286 520 290
rect 554 286 558 290
rect 1038 298 1042 302
rect 996 289 1000 296
rect 1054 289 1058 296
rect 1073 293 1077 297
rect 966 275 970 279
rect 189 266 193 270
rect 207 268 211 272
rect 267 268 271 272
rect 225 259 229 266
rect 283 259 287 266
rect 302 263 306 267
rect 320 268 324 272
rect 339 268 343 272
rect 399 268 403 272
rect 357 259 361 266
rect 415 259 419 266
rect 434 263 438 267
rect 452 268 456 272
rect 471 268 475 272
rect 531 268 535 272
rect 489 259 493 266
rect 1003 273 1007 277
rect 1023 273 1027 277
rect 1059 273 1063 277
rect 547 259 551 266
rect 568 263 572 267
rect 195 245 199 249
rect 232 243 236 247
rect 252 243 256 247
rect 288 243 292 247
rect 327 245 331 249
rect 364 243 368 247
rect 384 243 388 247
rect 420 243 424 247
rect 459 245 463 249
rect 496 243 500 247
rect 516 243 520 247
rect 552 243 556 247
rect 966 230 970 234
rect 1003 230 1007 234
rect 1023 230 1027 234
rect 1061 230 1065 234
rect 960 210 964 214
rect 978 212 982 216
rect 195 200 199 204
rect 232 200 236 204
rect 252 200 256 204
rect 290 200 294 204
rect 327 200 331 204
rect 364 200 368 204
rect 384 200 388 204
rect 422 200 426 204
rect 459 200 463 204
rect 496 200 500 204
rect 516 200 520 204
rect 554 200 558 204
rect 1038 212 1042 216
rect 996 203 1000 210
rect 1054 203 1058 210
rect 1073 207 1077 211
rect 1095 205 1099 209
rect 966 189 970 193
rect 189 180 193 184
rect 207 182 211 186
rect 267 182 271 186
rect 225 173 229 180
rect 283 173 287 180
rect 302 177 306 181
rect 320 182 324 186
rect 339 182 343 186
rect 399 182 403 186
rect 357 173 361 180
rect 415 173 419 180
rect 434 177 438 181
rect 452 182 456 186
rect 471 182 475 186
rect 531 182 535 186
rect 489 173 493 180
rect 1003 187 1007 191
rect 1023 187 1027 191
rect 1059 187 1063 191
rect 547 173 551 180
rect 568 177 572 181
rect 195 159 199 163
rect 232 157 236 161
rect 252 157 256 161
rect 288 157 292 161
rect 327 159 331 163
rect 364 157 368 161
rect 384 157 388 161
rect 420 157 424 161
rect 459 159 463 163
rect 496 157 500 161
rect 516 157 520 161
rect 552 157 556 161
rect 421 129 425 133
rect 445 129 449 133
rect 441 104 445 108
rect 456 96 460 100
rect 421 81 425 85
rect 445 81 449 85
rect 195 60 199 64
rect 232 60 236 64
rect 252 60 256 64
rect 290 60 294 64
rect 327 60 331 64
rect 364 60 368 64
rect 384 60 388 64
rect 422 60 426 64
rect 459 60 463 64
rect 496 60 500 64
rect 516 60 520 64
rect 554 60 558 64
rect 189 40 193 44
rect 207 42 211 46
rect 267 42 271 46
rect 225 33 229 40
rect 283 33 287 40
rect 302 37 306 41
rect 320 42 324 46
rect 339 42 343 46
rect 399 42 403 46
rect 357 33 361 40
rect 415 33 419 40
rect 434 37 438 41
rect 452 42 456 46
rect 471 42 475 46
rect 531 42 535 46
rect 489 33 493 40
rect 547 33 551 40
rect 568 37 572 41
rect 195 19 199 23
rect 232 17 236 21
rect 252 17 256 21
rect 288 17 292 21
rect 327 19 331 23
rect 364 17 368 21
rect 384 17 388 21
rect 420 17 424 21
rect 459 19 463 23
rect 496 17 500 21
rect 516 17 520 21
rect 552 17 556 21
<< metal1 >>
rect 648 975 663 979
rect 667 975 699 979
rect 703 975 766 979
rect 770 975 795 979
rect 799 975 831 979
rect 835 975 898 979
rect 902 975 927 979
rect 931 975 963 979
rect 967 975 1030 979
rect 1034 975 1059 979
rect 1063 975 1095 979
rect 1099 975 1162 979
rect 1166 975 1182 979
rect 588 968 687 972
rect 691 968 715 972
rect 719 968 745 972
rect 749 968 782 972
rect 786 968 819 972
rect 823 968 847 972
rect 851 968 877 972
rect 881 968 914 972
rect 918 968 951 972
rect 955 968 979 972
rect 983 968 1009 972
rect 1013 968 1046 972
rect 1050 968 1083 972
rect 1087 968 1111 972
rect 1115 968 1141 972
rect 1145 968 1178 972
rect 657 958 660 968
rect 678 958 681 968
rect 694 958 697 968
rect 708 961 713 965
rect 717 961 724 965
rect 736 958 739 968
rect 752 958 755 968
rect 773 958 776 968
rect 789 958 792 968
rect 810 958 813 968
rect 826 958 829 968
rect 840 961 845 965
rect 849 961 856 965
rect 868 958 871 968
rect 884 958 887 968
rect 905 958 908 968
rect 921 958 924 968
rect 942 958 945 968
rect 958 958 961 968
rect 972 961 977 965
rect 981 961 988 965
rect 1000 958 1003 968
rect 1016 958 1019 968
rect 1037 958 1040 968
rect 1053 958 1056 968
rect 1074 958 1077 968
rect 1090 958 1093 968
rect 1104 961 1109 965
rect 1113 961 1120 965
rect 1132 958 1135 968
rect 1148 958 1151 968
rect 1169 958 1172 968
rect 314 942 323 946
rect 327 942 359 946
rect 363 942 426 946
rect 430 942 642 946
rect 674 944 679 947
rect 683 944 707 947
rect 732 944 739 947
rect 743 944 765 947
rect 314 935 347 939
rect 351 935 375 939
rect 379 935 405 939
rect 409 935 442 939
rect 446 935 582 939
rect 317 925 320 935
rect 338 925 341 935
rect 354 925 357 935
rect 368 928 373 932
rect 377 928 384 932
rect 396 925 399 935
rect 412 925 415 935
rect 433 925 436 935
rect 690 934 697 937
rect 701 938 720 941
rect 720 931 723 937
rect 748 934 755 937
rect 759 938 776 941
rect 806 944 811 947
rect 815 944 839 947
rect 864 944 871 947
rect 875 944 897 947
rect 822 934 829 937
rect 833 938 852 941
rect 852 931 855 937
rect 880 934 887 937
rect 891 938 908 941
rect 938 944 943 947
rect 947 944 971 947
rect 996 944 1003 947
rect 1007 944 1029 947
rect 954 934 961 937
rect 965 938 984 941
rect 984 931 987 937
rect 1012 934 1019 937
rect 1023 938 1040 941
rect 1070 944 1075 947
rect 1079 944 1103 947
rect 1128 944 1135 947
rect 1139 944 1161 947
rect 1086 934 1093 937
rect 1097 938 1116 941
rect 312 908 321 912
rect 334 911 339 914
rect 343 911 367 914
rect 392 911 399 914
rect 403 911 425 914
rect 657 915 660 927
rect 678 915 681 927
rect 694 915 697 927
rect 708 918 720 921
rect 736 915 739 927
rect 752 915 755 927
rect 773 915 776 927
rect 789 915 792 927
rect 810 915 813 927
rect 826 915 829 927
rect 840 918 852 921
rect 868 915 871 927
rect 884 915 887 927
rect 905 915 908 927
rect 921 915 924 927
rect 942 915 945 927
rect 958 915 961 927
rect 972 918 984 921
rect 1000 915 1003 927
rect 1016 915 1019 927
rect 1037 915 1040 927
rect 1116 931 1119 937
rect 1144 934 1151 937
rect 1155 938 1172 941
rect 1053 915 1056 927
rect 1074 915 1077 927
rect 1090 915 1093 927
rect 1104 918 1116 921
rect 1132 915 1135 927
rect 1148 915 1151 927
rect 1169 915 1172 927
rect 600 911 687 915
rect 691 911 715 915
rect 719 911 745 915
rect 749 911 819 915
rect 823 911 847 915
rect 851 911 877 915
rect 881 911 951 915
rect 955 911 979 915
rect 983 911 1009 915
rect 1013 911 1083 915
rect 1087 911 1111 915
rect 1115 911 1141 915
rect 1145 911 1182 915
rect 350 901 357 904
rect 361 905 380 908
rect 380 898 383 904
rect 408 901 415 904
rect 419 905 434 908
rect 636 904 663 908
rect 667 904 714 908
rect 718 904 764 908
rect 768 904 795 908
rect 799 904 846 908
rect 850 904 896 908
rect 900 904 927 908
rect 931 904 978 908
rect 982 904 1028 908
rect 1032 904 1059 908
rect 1063 904 1110 908
rect 1114 904 1160 908
rect 1164 904 1182 908
rect 317 882 320 894
rect 338 882 341 894
rect 354 882 357 894
rect 368 885 380 888
rect 396 882 399 894
rect 412 882 415 894
rect 433 882 436 894
rect 588 891 661 895
rect 665 891 677 895
rect 681 891 695 895
rect 699 891 706 895
rect 710 891 712 895
rect 716 891 731 895
rect 735 891 768 895
rect 772 891 773 895
rect 777 891 785 895
rect 789 891 813 895
rect 817 891 829 895
rect 833 891 853 895
rect 857 891 907 895
rect 911 891 934 895
rect 938 891 988 895
rect 992 891 1011 895
rect 624 884 688 888
rect 692 884 719 888
rect 723 884 741 888
rect 745 884 806 888
rect 810 884 824 888
rect 836 887 839 891
rect 314 878 347 882
rect 351 878 375 882
rect 379 878 405 882
rect 409 878 594 882
rect 314 871 323 875
rect 327 871 374 875
rect 378 871 424 875
rect 428 871 630 875
rect 731 877 734 881
rect 758 877 759 881
rect 803 877 805 881
rect 845 874 848 879
rect 860 881 863 891
rect 890 887 893 891
rect 917 887 920 891
rect 312 855 328 859
rect 437 857 441 861
rect 453 857 457 861
rect 461 857 663 861
rect 671 860 674 866
rect 678 860 681 866
rect 671 857 681 860
rect 671 852 674 857
rect 320 848 324 852
rect 336 848 457 852
rect 678 852 681 857
rect 687 862 690 866
rect 687 858 689 862
rect 693 858 695 862
rect 703 861 706 866
rect 731 863 734 866
rect 703 859 714 861
rect 687 852 690 858
rect 703 857 709 859
rect 703 852 706 857
rect 713 857 714 859
rect 732 859 734 863
rect 731 852 734 859
rect 834 870 837 873
rect 876 870 879 873
rect 747 862 750 866
rect 757 862 760 866
rect 757 858 766 862
rect 778 861 781 866
rect 803 862 806 866
rect 747 852 750 858
rect 757 852 760 858
rect 778 857 779 861
rect 783 857 786 860
rect 805 858 806 862
rect 821 861 824 866
rect 845 865 848 870
rect 853 866 864 869
rect 876 867 884 870
rect 778 852 781 857
rect 803 852 806 858
rect 821 852 824 857
rect 307 840 323 844
rect 327 840 390 844
rect 394 840 426 844
rect 430 840 642 844
rect 723 839 724 843
rect 748 840 749 844
rect 795 839 796 843
rect 311 833 344 837
rect 348 833 374 837
rect 378 833 402 837
rect 406 833 582 837
rect 317 823 320 833
rect 338 823 341 833
rect 354 823 357 833
rect 369 826 376 830
rect 380 826 385 830
rect 396 823 399 833
rect 412 823 415 833
rect 433 823 436 833
rect 612 832 676 836
rect 680 832 735 836
rect 739 832 760 836
rect 764 832 791 836
rect 795 832 824 836
rect 836 829 839 861
rect 853 860 856 866
rect 876 861 879 867
rect 888 862 891 865
rect 899 865 902 879
rect 926 874 929 879
rect 941 881 944 891
rect 971 887 974 891
rect 910 870 911 873
rect 915 870 918 873
rect 957 870 960 873
rect 899 862 907 865
rect 926 865 929 870
rect 899 857 902 862
rect 907 858 911 862
rect 934 866 945 869
rect 957 867 965 870
rect 851 851 856 856
rect 860 829 863 857
rect 890 829 893 853
rect 917 829 920 861
rect 934 860 937 866
rect 957 861 960 867
rect 969 862 972 865
rect 980 865 983 879
rect 980 862 992 865
rect 980 857 983 862
rect 932 851 937 856
rect 941 829 944 857
rect 971 829 974 853
rect 600 825 662 829
rect 666 825 668 829
rect 672 825 676 829
rect 680 825 694 829
rect 698 825 703 829
rect 707 825 712 829
rect 716 825 735 829
rect 739 825 769 829
rect 773 825 784 829
rect 788 825 812 829
rect 816 825 829 829
rect 833 825 853 829
rect 857 825 907 829
rect 914 825 934 829
rect 938 825 988 829
rect 328 809 350 812
rect 354 809 361 812
rect 612 818 676 822
rect 680 818 735 822
rect 739 818 760 822
rect 764 818 791 822
rect 795 818 824 822
rect 386 809 410 812
rect 414 809 419 812
rect 723 811 724 815
rect 748 810 749 814
rect 795 811 796 815
rect 432 806 441 810
rect 319 803 334 806
rect 373 803 392 806
rect 338 799 345 802
rect 370 796 373 802
rect 396 799 403 802
rect 671 797 674 802
rect 678 797 681 802
rect 661 794 663 797
rect 671 794 681 797
rect 317 780 320 792
rect 338 780 341 792
rect 354 780 357 792
rect 373 783 385 786
rect 396 780 399 792
rect 412 780 415 792
rect 433 780 436 792
rect 671 788 674 794
rect 678 788 681 794
rect 687 796 690 802
rect 703 797 706 802
rect 687 792 689 796
rect 693 792 695 796
rect 703 795 709 797
rect 713 795 714 797
rect 703 793 714 795
rect 731 795 734 802
rect 687 788 690 792
rect 703 788 706 793
rect 732 791 734 795
rect 731 788 734 791
rect 747 796 750 802
rect 757 796 760 802
rect 778 797 781 802
rect 757 792 766 796
rect 778 793 779 797
rect 783 794 786 797
rect 803 796 806 802
rect 821 797 824 802
rect 860 805 863 825
rect 941 805 944 825
rect 747 788 750 792
rect 757 788 760 792
rect 778 788 781 793
rect 805 792 806 796
rect 803 788 806 792
rect 821 788 824 793
rect 851 792 856 797
rect 860 793 861 796
rect 876 795 879 801
rect 876 792 884 795
rect 931 792 936 797
rect 940 793 942 796
rect 957 795 960 801
rect 957 792 965 795
rect 876 789 879 792
rect 957 789 960 792
rect 307 776 344 780
rect 348 776 374 780
rect 378 776 402 780
rect 406 776 594 780
rect 731 773 734 777
rect 758 773 759 777
rect 803 773 805 777
rect 307 769 325 773
rect 329 769 375 773
rect 379 769 426 773
rect 430 769 630 773
rect 676 766 688 770
rect 692 766 719 770
rect 723 766 741 770
rect 745 766 806 770
rect 810 766 824 770
rect 860 763 863 781
rect 941 763 944 781
rect 588 759 661 763
rect 665 759 677 763
rect 681 759 695 763
rect 699 759 706 763
rect 710 759 712 763
rect 716 759 731 763
rect 735 759 768 763
rect 772 759 773 763
rect 777 759 785 763
rect 789 759 813 763
rect 817 759 829 763
rect 833 759 853 763
rect 857 759 907 763
rect 911 759 934 763
rect 938 759 996 763
rect 1000 759 1011 763
rect 624 752 672 756
rect 676 752 688 756
rect 692 752 719 756
rect 723 752 741 756
rect 745 752 806 756
rect 810 752 824 756
rect 860 749 863 759
rect 890 755 893 759
rect 941 755 944 759
rect 731 745 734 749
rect 758 745 759 749
rect 803 745 805 749
rect 660 725 663 728
rect 671 728 674 734
rect 678 728 681 734
rect 671 725 681 728
rect 671 720 674 725
rect 678 720 681 725
rect 687 730 690 734
rect 687 726 689 730
rect 693 726 695 730
rect 703 729 706 734
rect 731 731 734 734
rect 703 727 714 729
rect 687 720 690 726
rect 703 725 709 727
rect 703 720 706 725
rect 713 725 714 727
rect 732 727 734 731
rect 731 720 734 727
rect 876 738 879 741
rect 747 730 750 734
rect 757 730 760 734
rect 757 726 766 730
rect 778 729 781 734
rect 803 730 806 734
rect 747 720 750 726
rect 757 720 760 726
rect 778 725 779 729
rect 783 725 786 728
rect 805 726 806 730
rect 821 729 824 734
rect 853 734 864 737
rect 876 735 884 738
rect 778 720 781 725
rect 803 720 806 726
rect 853 728 856 734
rect 876 729 879 735
rect 888 730 891 733
rect 899 733 902 747
rect 950 742 953 747
rect 965 749 968 759
rect 995 755 998 759
rect 934 738 935 741
rect 939 738 942 741
rect 981 738 984 741
rect 907 733 912 738
rect 950 733 953 738
rect 899 730 907 733
rect 821 720 824 725
rect 899 725 902 730
rect 958 734 969 737
rect 981 735 989 738
rect 851 719 856 724
rect 723 707 724 711
rect 748 708 749 712
rect 795 707 796 711
rect 612 700 676 704
rect 680 700 735 704
rect 739 700 760 704
rect 764 700 791 704
rect 795 700 824 704
rect 860 697 863 725
rect 890 697 893 721
rect 941 697 944 729
rect 958 728 961 734
rect 981 729 984 735
rect 993 730 996 733
rect 1004 733 1007 747
rect 1004 730 1010 733
rect 1004 725 1007 730
rect 956 719 961 724
rect 965 697 968 725
rect 995 697 998 721
rect 600 693 662 697
rect 666 693 668 697
rect 672 693 676 697
rect 680 693 694 697
rect 698 693 703 697
rect 707 693 712 697
rect 716 693 735 697
rect 739 693 769 697
rect 773 693 784 697
rect 788 693 812 697
rect 816 693 829 697
rect 833 693 853 697
rect 857 693 907 697
rect 911 693 934 697
rect 938 693 958 697
rect 962 693 1010 697
rect 612 686 676 690
rect 680 686 735 690
rect 739 686 760 690
rect 764 686 791 690
rect 795 686 824 690
rect 723 679 724 683
rect 748 678 749 682
rect 795 679 796 683
rect 860 674 863 693
rect 965 674 968 693
rect 671 665 674 670
rect 678 665 681 670
rect 661 662 663 665
rect 671 662 681 665
rect 671 656 674 662
rect 678 656 681 662
rect 687 664 690 670
rect 703 665 706 670
rect 687 660 689 664
rect 693 660 695 664
rect 703 663 709 665
rect 713 663 714 665
rect 703 661 714 663
rect 731 663 734 670
rect 687 656 690 660
rect 703 656 706 661
rect 732 659 734 663
rect 731 656 734 659
rect 747 664 750 670
rect 757 664 760 670
rect 778 665 781 670
rect 757 660 766 664
rect 778 661 779 665
rect 783 662 786 665
rect 803 664 806 670
rect 821 665 824 670
rect 747 656 750 660
rect 757 656 760 660
rect 778 656 781 661
rect 805 660 806 664
rect 850 661 855 666
rect 859 662 861 665
rect 876 664 879 670
rect 876 661 884 664
rect 956 661 961 666
rect 965 662 966 665
rect 981 664 984 670
rect 981 661 989 664
rect 803 656 806 660
rect 821 656 824 661
rect 876 658 879 661
rect 981 658 984 661
rect 731 641 734 645
rect 758 641 759 645
rect 803 641 805 645
rect 624 634 688 638
rect 692 634 719 638
rect 723 634 741 638
rect 745 634 806 638
rect 810 634 824 638
rect 860 631 863 650
rect 965 631 968 650
rect 588 627 661 631
rect 665 627 677 631
rect 681 627 695 631
rect 699 627 706 631
rect 710 627 712 631
rect 716 627 731 631
rect 735 627 768 631
rect 772 627 773 631
rect 777 627 785 631
rect 789 627 813 631
rect 817 627 829 631
rect 833 627 853 631
rect 857 627 907 631
rect 911 627 934 631
rect 938 627 988 631
rect 992 627 996 631
rect 1000 627 1024 631
rect 1028 627 1078 631
rect 624 620 688 624
rect 692 620 719 624
rect 723 620 741 624
rect 745 620 806 624
rect 810 620 824 624
rect 860 617 863 627
rect 890 623 893 627
rect 917 623 920 627
rect 731 613 734 617
rect 758 613 759 617
rect 803 613 805 617
rect 660 593 663 596
rect 671 596 674 602
rect 678 596 681 602
rect 671 593 681 596
rect 671 588 674 593
rect 678 588 681 593
rect 687 598 690 602
rect 687 594 689 598
rect 693 594 695 598
rect 703 597 706 602
rect 731 599 734 602
rect 703 595 714 597
rect 687 588 690 594
rect 703 593 709 595
rect 703 588 706 593
rect 713 593 714 595
rect 732 595 734 599
rect 731 588 734 595
rect 876 606 879 609
rect 747 598 750 602
rect 757 598 760 602
rect 757 594 766 598
rect 778 597 781 602
rect 803 598 806 602
rect 747 588 750 594
rect 757 588 760 594
rect 778 593 779 597
rect 783 593 786 596
rect 805 594 806 598
rect 821 597 824 602
rect 853 602 864 605
rect 876 603 884 606
rect 778 588 781 593
rect 803 588 806 594
rect 853 596 856 602
rect 876 597 879 603
rect 888 598 891 601
rect 899 601 902 615
rect 926 610 929 615
rect 941 617 944 627
rect 971 623 974 627
rect 1007 623 1010 627
rect 910 606 911 609
rect 915 606 918 609
rect 957 606 960 609
rect 899 598 907 601
rect 926 601 929 606
rect 821 588 824 593
rect 899 593 902 598
rect 907 594 911 598
rect 934 602 945 605
rect 957 603 965 606
rect 851 587 856 592
rect 723 575 724 579
rect 748 576 749 580
rect 795 575 796 579
rect 612 568 676 572
rect 680 568 735 572
rect 739 568 760 572
rect 764 568 791 572
rect 795 568 824 572
rect 860 565 863 593
rect 890 565 893 589
rect 917 565 920 597
rect 934 596 937 602
rect 957 597 960 603
rect 969 598 972 601
rect 980 601 983 615
rect 1016 610 1019 615
rect 1031 617 1034 627
rect 1061 623 1064 627
rect 1005 606 1008 609
rect 1047 606 1050 609
rect 980 598 989 601
rect 1016 601 1019 606
rect 980 593 983 598
rect 932 587 937 592
rect 941 565 944 593
rect 1023 604 1035 605
rect 1027 602 1035 604
rect 1047 603 1055 606
rect 1047 597 1050 603
rect 1059 598 1062 601
rect 1070 601 1073 615
rect 1070 598 1090 601
rect 971 565 974 589
rect 1007 565 1010 597
rect 1070 593 1073 598
rect 1031 565 1034 593
rect 1061 565 1064 589
rect 600 561 662 565
rect 666 561 668 565
rect 672 561 676 565
rect 680 561 694 565
rect 698 561 703 565
rect 707 561 712 565
rect 716 561 735 565
rect 739 561 769 565
rect 773 561 784 565
rect 788 561 812 565
rect 816 561 829 565
rect 833 561 853 565
rect 857 561 907 565
rect 914 561 934 565
rect 938 561 988 565
rect 992 561 1024 565
rect 1028 561 1078 565
rect 612 554 676 558
rect 680 554 735 558
rect 739 554 760 558
rect 764 554 791 558
rect 795 554 824 558
rect 723 547 724 551
rect 748 546 749 550
rect 795 547 796 551
rect 671 533 674 538
rect 678 533 681 538
rect 661 530 663 533
rect 671 530 681 533
rect 671 524 674 530
rect 678 524 681 530
rect 687 532 690 538
rect 703 533 706 538
rect 687 528 689 532
rect 693 528 695 532
rect 703 531 709 533
rect 713 531 714 533
rect 703 529 714 531
rect 731 531 734 538
rect 687 524 690 528
rect 703 524 706 529
rect 732 527 734 531
rect 731 524 734 527
rect 747 532 750 538
rect 757 532 760 538
rect 778 533 781 538
rect 757 528 766 532
rect 778 529 779 533
rect 783 530 786 533
rect 803 532 806 538
rect 821 533 824 538
rect 860 539 863 561
rect 941 539 944 561
rect 1031 539 1034 561
rect 747 524 750 528
rect 757 524 760 528
rect 778 524 781 529
rect 805 528 806 532
rect 803 524 806 528
rect 821 524 824 529
rect 851 526 856 531
rect 860 527 861 530
rect 876 529 879 535
rect 876 526 884 529
rect 931 526 936 531
rect 940 527 942 530
rect 957 529 960 535
rect 957 526 965 529
rect 1024 527 1032 530
rect 1047 529 1050 535
rect 1047 526 1055 529
rect 876 523 879 526
rect 957 523 960 526
rect 1047 523 1050 526
rect 731 509 734 513
rect 758 509 759 513
rect 803 509 805 513
rect 624 502 688 506
rect 692 502 719 506
rect 723 502 741 506
rect 745 502 806 506
rect 810 502 824 506
rect 860 499 863 515
rect 941 499 944 515
rect 1031 499 1034 515
rect 588 495 661 499
rect 665 495 677 499
rect 681 495 695 499
rect 699 495 706 499
rect 710 495 712 499
rect 716 495 731 499
rect 735 495 768 499
rect 772 495 773 499
rect 777 495 785 499
rect 789 495 813 499
rect 817 495 829 499
rect 833 495 853 499
rect 857 495 907 499
rect 911 495 934 499
rect 938 495 1024 499
rect 1028 495 1082 499
rect 624 488 688 492
rect 692 488 719 492
rect 723 488 741 492
rect 745 488 806 492
rect 810 488 824 492
rect 860 485 863 495
rect 890 491 893 495
rect 731 481 734 485
rect 758 481 759 485
rect 803 481 805 485
rect 660 461 663 464
rect 671 464 674 470
rect 678 464 681 470
rect 671 461 681 464
rect 671 456 674 461
rect 678 456 681 461
rect 687 466 690 470
rect 687 462 689 466
rect 693 462 695 466
rect 703 465 706 470
rect 731 467 734 470
rect 703 463 714 465
rect 687 456 690 462
rect 703 461 709 463
rect 703 456 706 461
rect 713 461 714 463
rect 732 463 734 467
rect 731 456 734 463
rect 876 474 879 477
rect 747 466 750 470
rect 757 466 760 470
rect 757 462 766 466
rect 778 465 781 470
rect 803 466 806 470
rect 747 456 750 462
rect 757 456 760 462
rect 778 461 779 465
rect 783 461 786 464
rect 805 462 806 466
rect 821 465 824 470
rect 853 470 864 473
rect 876 471 884 474
rect 778 456 781 461
rect 803 456 806 462
rect 853 464 856 470
rect 876 465 879 471
rect 888 466 891 469
rect 899 469 902 483
rect 907 469 912 474
rect 899 466 907 469
rect 821 456 824 461
rect 899 461 902 466
rect 851 455 856 460
rect 182 440 191 444
rect 195 440 227 444
rect 231 440 294 444
rect 298 440 323 444
rect 327 440 359 444
rect 363 440 426 444
rect 430 440 455 444
rect 459 440 491 444
rect 495 440 558 444
rect 562 440 642 444
rect 723 443 724 447
rect 748 444 749 448
rect 795 443 796 447
rect 182 433 215 437
rect 219 433 243 437
rect 247 433 273 437
rect 277 433 310 437
rect 314 433 347 437
rect 351 433 375 437
rect 379 433 405 437
rect 409 433 442 437
rect 446 433 479 437
rect 483 433 507 437
rect 511 433 537 437
rect 541 433 574 437
rect 578 433 582 437
rect 655 436 676 440
rect 680 436 685 440
rect 689 436 735 440
rect 739 436 760 440
rect 764 436 791 440
rect 795 436 824 440
rect 860 433 863 461
rect 890 433 893 457
rect 185 423 188 433
rect 206 423 209 433
rect 222 423 225 433
rect 236 426 241 430
rect 245 426 252 430
rect 264 423 267 433
rect 280 423 283 433
rect 301 423 304 433
rect 317 423 320 433
rect 338 423 341 433
rect 354 423 357 433
rect 368 426 373 430
rect 377 426 384 430
rect 396 423 399 433
rect 412 423 415 433
rect 433 423 436 433
rect 449 423 452 433
rect 470 423 473 433
rect 486 423 489 433
rect 500 426 505 430
rect 509 426 516 430
rect 528 423 531 433
rect 544 423 547 433
rect 565 423 568 433
rect 600 429 662 433
rect 666 429 668 433
rect 672 429 676 433
rect 680 429 694 433
rect 698 429 703 433
rect 707 429 712 433
rect 716 429 735 433
rect 739 429 769 433
rect 773 429 784 433
rect 788 429 812 433
rect 816 429 829 433
rect 833 429 853 433
rect 857 429 937 433
rect 941 429 955 433
rect 959 429 964 433
rect 968 429 973 433
rect 977 429 996 433
rect 1000 429 1030 433
rect 1034 429 1045 433
rect 1049 429 1073 433
rect 1077 429 1086 433
rect 202 409 207 412
rect 211 409 235 412
rect 260 409 267 412
rect 271 409 293 412
rect 313 409 320 412
rect 334 409 339 412
rect 343 409 367 412
rect 392 409 399 412
rect 403 409 425 412
rect 445 409 452 412
rect 466 409 471 412
rect 475 409 499 412
rect 612 422 676 426
rect 680 422 685 426
rect 689 422 735 426
rect 739 422 760 426
rect 764 422 791 426
rect 795 422 824 426
rect 524 409 531 412
rect 535 409 557 412
rect 723 415 724 419
rect 748 414 749 418
rect 795 415 796 419
rect 218 399 225 402
rect 229 403 248 406
rect 248 396 251 402
rect 276 399 283 402
rect 287 403 302 406
rect 350 399 357 402
rect 361 403 380 406
rect 380 396 383 402
rect 408 399 415 402
rect 419 403 434 406
rect 482 399 489 402
rect 493 403 512 406
rect 512 396 515 402
rect 540 399 547 402
rect 551 403 568 406
rect 671 401 674 406
rect 678 401 681 406
rect 661 398 663 401
rect 671 398 681 401
rect 671 392 674 398
rect 185 380 188 392
rect 206 380 209 392
rect 222 380 225 392
rect 236 383 248 386
rect 264 380 267 392
rect 280 380 283 392
rect 301 380 304 392
rect 317 380 320 392
rect 338 380 341 392
rect 354 380 357 392
rect 368 383 380 386
rect 396 380 399 392
rect 412 380 415 392
rect 433 380 436 392
rect 449 380 452 392
rect 470 380 473 392
rect 486 380 489 392
rect 500 383 512 386
rect 528 380 531 392
rect 544 380 547 392
rect 565 380 568 392
rect 678 392 681 398
rect 687 400 690 406
rect 703 401 706 406
rect 687 396 689 400
rect 693 396 695 400
rect 703 399 709 401
rect 713 399 714 401
rect 703 397 714 399
rect 731 399 734 406
rect 687 392 690 396
rect 703 392 706 397
rect 732 395 734 399
rect 731 392 734 395
rect 747 400 750 406
rect 757 400 760 406
rect 778 401 781 406
rect 757 396 766 400
rect 778 397 779 401
rect 783 398 786 401
rect 803 400 806 406
rect 821 401 824 406
rect 860 403 863 429
rect 896 422 915 426
rect 919 422 937 426
rect 941 422 996 426
rect 1000 422 1021 426
rect 1025 422 1052 426
rect 1056 422 1085 426
rect 896 410 899 422
rect 984 415 985 419
rect 1009 414 1010 418
rect 1056 415 1057 419
rect 747 392 750 396
rect 757 392 760 396
rect 778 392 781 397
rect 805 396 806 400
rect 923 401 926 406
rect 932 401 935 406
rect 939 401 942 406
rect 803 392 806 396
rect 821 392 824 397
rect 850 390 855 395
rect 859 391 861 394
rect 876 393 879 399
rect 908 398 942 401
rect 876 390 884 393
rect 876 387 879 390
rect 182 376 215 380
rect 219 376 243 380
rect 247 376 273 380
rect 277 376 347 380
rect 351 376 375 380
rect 379 376 405 380
rect 409 376 479 380
rect 483 376 507 380
rect 511 376 537 380
rect 541 376 594 380
rect 731 377 734 381
rect 758 377 759 381
rect 803 377 805 381
rect 908 384 911 398
rect 932 392 935 398
rect 939 392 942 398
rect 948 400 951 406
rect 964 401 967 406
rect 948 396 950 400
rect 954 396 956 400
rect 964 399 970 401
rect 974 399 975 401
rect 964 397 975 399
rect 992 399 995 406
rect 948 392 951 396
rect 964 392 967 397
rect 993 395 995 399
rect 992 392 995 395
rect 1008 400 1011 406
rect 1018 400 1021 406
rect 1039 401 1042 406
rect 1018 396 1027 400
rect 1039 397 1040 401
rect 1044 398 1047 401
rect 1064 400 1067 406
rect 1082 401 1085 406
rect 1008 392 1011 396
rect 1018 392 1021 396
rect 1039 392 1042 397
rect 1066 396 1067 400
rect 1064 392 1067 396
rect 1082 392 1085 397
rect 182 369 191 373
rect 195 369 242 373
rect 246 369 292 373
rect 296 369 323 373
rect 327 369 374 373
rect 378 369 424 373
rect 428 369 455 373
rect 459 369 506 373
rect 510 369 556 373
rect 560 370 630 373
rect 674 370 688 374
rect 692 370 719 374
rect 723 370 741 374
rect 745 370 806 374
rect 810 370 824 374
rect 860 367 863 379
rect 992 377 995 381
rect 1019 377 1020 381
rect 1064 377 1066 381
rect 900 370 905 374
rect 909 370 949 374
rect 953 370 980 374
rect 984 370 1002 374
rect 1006 370 1067 374
rect 1071 370 1085 374
rect 189 363 573 366
rect 588 363 661 367
rect 665 363 677 367
rect 681 363 695 367
rect 699 363 706 367
rect 710 363 712 367
rect 716 363 731 367
rect 735 363 768 367
rect 772 363 773 367
rect 777 363 785 367
rect 789 363 813 367
rect 817 363 853 367
rect 857 363 896 367
rect 900 363 907 367
rect 911 363 922 367
rect 926 363 938 367
rect 942 363 956 367
rect 960 363 967 367
rect 971 363 973 367
rect 977 363 992 367
rect 996 363 1029 367
rect 1033 363 1034 367
rect 1038 363 1046 367
rect 1050 363 1074 367
rect 1078 363 1086 367
rect 332 356 441 359
rect 624 356 670 360
rect 674 356 904 359
rect 1094 357 1102 361
rect 312 348 316 352
rect 320 348 324 352
rect 612 349 914 352
rect 1090 341 1094 345
rect 172 337 300 341
rect 304 337 320 341
rect 336 337 1115 341
rect 328 330 573 333
rect 648 330 962 334
rect 966 330 998 334
rect 1002 330 1065 334
rect 1069 330 1085 334
rect 343 323 573 326
rect 588 323 948 327
rect 952 323 986 327
rect 990 323 1014 327
rect 1018 323 1044 327
rect 1048 323 1081 327
rect 312 314 316 318
rect 320 314 324 318
rect 956 313 959 323
rect 977 313 980 323
rect 993 313 996 323
rect 1007 316 1012 320
rect 1016 316 1023 320
rect 1035 313 1038 323
rect 1051 313 1054 323
rect 1072 313 1075 323
rect 332 307 442 310
rect 182 300 191 304
rect 195 300 227 304
rect 231 300 294 304
rect 298 300 323 304
rect 327 300 359 304
rect 363 300 426 304
rect 430 300 455 304
rect 459 300 491 304
rect 495 300 558 304
rect 562 300 642 304
rect 182 293 215 297
rect 219 293 243 297
rect 247 293 273 297
rect 277 293 310 297
rect 314 293 347 297
rect 351 293 375 297
rect 379 293 405 297
rect 409 293 442 297
rect 446 293 479 297
rect 483 293 507 297
rect 511 293 537 297
rect 541 293 574 297
rect 578 293 582 297
rect 973 299 978 302
rect 982 299 1006 302
rect 1031 299 1038 302
rect 1042 299 1064 302
rect 185 283 188 293
rect 206 283 209 293
rect 222 283 225 293
rect 236 286 241 290
rect 245 286 252 290
rect 264 283 267 293
rect 280 283 283 293
rect 301 283 304 293
rect 317 283 320 293
rect 338 283 341 293
rect 354 283 357 293
rect 368 286 373 290
rect 377 286 384 290
rect 396 283 399 293
rect 412 283 415 293
rect 433 283 436 293
rect 449 283 452 293
rect 470 283 473 293
rect 486 283 489 293
rect 500 286 505 290
rect 509 286 516 290
rect 528 283 531 293
rect 544 283 547 293
rect 565 283 568 293
rect 989 289 996 292
rect 1000 293 1019 296
rect 202 269 207 272
rect 211 269 235 272
rect 260 269 267 272
rect 271 269 293 272
rect 313 269 320 272
rect 334 269 339 272
rect 343 269 367 272
rect 392 269 399 272
rect 403 269 425 272
rect 445 269 452 272
rect 466 269 471 272
rect 475 269 499 272
rect 524 269 531 272
rect 535 269 557 272
rect 1019 286 1022 292
rect 1047 289 1054 292
rect 1058 293 1073 296
rect 956 270 959 282
rect 977 270 980 282
rect 993 270 996 282
rect 1007 273 1019 276
rect 1035 270 1038 282
rect 1051 270 1054 282
rect 1072 270 1075 282
rect 218 259 225 262
rect 229 263 248 266
rect 248 256 251 262
rect 276 259 283 262
rect 287 263 302 266
rect 350 259 357 262
rect 361 263 380 266
rect 380 256 383 262
rect 408 259 415 262
rect 419 263 434 266
rect 482 259 489 262
rect 493 263 512 266
rect 512 256 515 262
rect 540 259 547 262
rect 551 263 568 266
rect 600 266 986 270
rect 990 266 1014 270
rect 1018 266 1044 270
rect 1048 266 1085 270
rect 636 259 962 263
rect 966 259 1013 263
rect 1017 259 1063 263
rect 1067 259 1085 263
rect 185 240 188 252
rect 206 240 209 252
rect 222 240 225 252
rect 236 243 248 246
rect 264 240 267 252
rect 280 240 283 252
rect 301 240 304 252
rect 317 240 320 252
rect 338 240 341 252
rect 354 240 357 252
rect 368 243 380 246
rect 396 240 399 252
rect 412 240 415 252
rect 433 240 436 252
rect 449 240 452 252
rect 470 240 473 252
rect 486 240 489 252
rect 500 243 512 246
rect 528 240 531 252
rect 544 240 547 252
rect 565 240 568 252
rect 959 252 1080 255
rect 648 244 962 248
rect 966 244 998 248
rect 1002 244 1065 248
rect 1069 244 1085 248
rect 182 236 215 240
rect 219 236 243 240
rect 247 236 273 240
rect 277 236 347 240
rect 351 236 375 240
rect 379 236 405 240
rect 409 236 479 240
rect 483 236 507 240
rect 511 236 537 240
rect 541 236 594 240
rect 952 237 986 241
rect 990 237 1014 241
rect 1018 237 1044 241
rect 1048 237 1081 241
rect 182 229 191 233
rect 195 229 242 233
rect 246 229 292 233
rect 296 229 323 233
rect 327 229 374 233
rect 378 229 424 233
rect 428 229 455 233
rect 459 229 506 233
rect 510 229 556 233
rect 560 229 630 233
rect 956 227 959 237
rect 977 227 980 237
rect 993 227 996 237
rect 1007 230 1012 234
rect 1016 230 1023 234
rect 1035 227 1038 237
rect 1051 227 1054 237
rect 1072 227 1075 237
rect 188 222 573 225
rect 182 214 191 218
rect 195 214 227 218
rect 231 214 294 218
rect 298 214 323 218
rect 327 214 359 218
rect 363 214 426 218
rect 430 214 455 218
rect 459 214 491 218
rect 495 214 558 218
rect 562 214 642 218
rect 182 207 215 211
rect 219 207 243 211
rect 247 207 273 211
rect 277 207 310 211
rect 314 207 347 211
rect 351 207 375 211
rect 379 207 405 211
rect 409 207 442 211
rect 446 207 479 211
rect 483 207 507 211
rect 511 207 537 211
rect 541 207 574 211
rect 578 207 582 211
rect 973 213 978 216
rect 982 213 1006 216
rect 1031 213 1038 216
rect 1042 213 1064 216
rect 185 197 188 207
rect 206 197 209 207
rect 222 197 225 207
rect 236 200 241 204
rect 245 200 252 204
rect 264 197 267 207
rect 280 197 283 207
rect 301 197 304 207
rect 317 197 320 207
rect 338 197 341 207
rect 354 197 357 207
rect 368 200 373 204
rect 377 200 384 204
rect 396 197 399 207
rect 412 197 415 207
rect 433 197 436 207
rect 449 197 452 207
rect 470 197 473 207
rect 486 197 489 207
rect 500 200 505 204
rect 509 200 516 204
rect 528 197 531 207
rect 544 197 547 207
rect 565 197 568 207
rect 989 203 996 206
rect 1000 207 1019 210
rect 202 183 207 186
rect 211 183 235 186
rect 260 183 267 186
rect 271 183 293 186
rect 313 183 320 186
rect 334 183 339 186
rect 343 183 367 186
rect 392 183 399 186
rect 403 183 425 186
rect 445 183 452 186
rect 466 183 471 186
rect 475 183 499 186
rect 524 183 531 186
rect 535 183 557 186
rect 1019 200 1022 206
rect 1047 203 1054 206
rect 1058 207 1073 210
rect 1084 205 1095 209
rect 956 184 959 196
rect 977 184 980 196
rect 993 184 996 196
rect 1007 187 1019 190
rect 1035 184 1038 196
rect 1051 184 1054 196
rect 1072 184 1075 196
rect 218 173 225 176
rect 229 177 248 180
rect 248 170 251 176
rect 276 173 283 176
rect 287 177 302 180
rect 350 173 357 176
rect 361 177 380 180
rect 380 170 383 176
rect 408 173 415 176
rect 419 177 434 180
rect 482 173 489 176
rect 493 177 512 180
rect 512 170 515 176
rect 540 173 547 176
rect 551 177 568 180
rect 600 180 986 184
rect 990 180 1014 184
rect 1018 180 1044 184
rect 1048 180 1085 184
rect 636 173 962 177
rect 966 173 1013 177
rect 1017 173 1063 177
rect 1067 173 1085 177
rect 185 154 188 166
rect 206 154 209 166
rect 222 154 225 166
rect 236 157 248 160
rect 264 154 267 166
rect 280 154 283 166
rect 301 154 304 166
rect 317 154 320 166
rect 338 154 341 166
rect 354 154 357 166
rect 368 157 380 160
rect 396 154 399 166
rect 412 154 415 166
rect 433 154 436 166
rect 449 154 452 166
rect 470 154 473 166
rect 486 154 489 166
rect 500 157 512 160
rect 528 154 531 166
rect 544 154 547 166
rect 565 154 568 166
rect 182 150 215 154
rect 219 150 243 154
rect 247 150 273 154
rect 277 150 347 154
rect 351 150 375 154
rect 379 150 405 154
rect 409 150 479 154
rect 483 150 507 154
rect 511 150 537 154
rect 541 150 594 154
rect 182 143 191 147
rect 195 143 242 147
rect 246 143 292 147
rect 296 143 323 147
rect 327 143 374 147
rect 378 143 424 147
rect 428 143 455 147
rect 459 143 506 147
rect 510 143 556 147
rect 560 143 630 147
rect 188 137 573 140
rect 313 130 417 133
rect 429 122 433 126
rect 437 122 441 126
rect 172 111 417 115
rect 421 111 437 115
rect 453 111 1102 115
rect 1106 111 1115 115
rect 445 104 573 107
rect 460 97 573 100
rect 429 88 433 92
rect 437 88 441 92
rect 313 81 417 84
rect 182 74 191 78
rect 195 74 227 78
rect 231 74 294 78
rect 298 74 323 78
rect 327 74 359 78
rect 363 74 426 78
rect 430 74 455 78
rect 459 74 491 78
rect 495 74 558 78
rect 562 74 642 78
rect 182 67 215 71
rect 219 67 243 71
rect 247 67 273 71
rect 277 67 310 71
rect 314 67 347 71
rect 351 67 375 71
rect 379 67 405 71
rect 409 67 442 71
rect 446 67 479 71
rect 483 67 507 71
rect 511 67 537 71
rect 541 67 574 71
rect 578 67 582 71
rect 185 57 188 67
rect 206 57 209 67
rect 222 57 225 67
rect 236 60 241 64
rect 245 60 252 64
rect 264 57 267 67
rect 280 57 283 67
rect 301 57 304 67
rect 317 57 320 67
rect 338 57 341 67
rect 354 57 357 67
rect 368 60 373 64
rect 377 60 384 64
rect 396 57 399 67
rect 412 57 415 67
rect 433 57 436 67
rect 449 57 452 67
rect 470 57 473 67
rect 486 57 489 67
rect 500 60 505 64
rect 509 60 516 64
rect 528 57 531 67
rect 544 57 547 67
rect 565 57 568 67
rect 202 43 207 46
rect 211 43 235 46
rect 260 43 267 46
rect 271 43 293 46
rect 313 43 320 46
rect 334 43 339 46
rect 343 43 367 46
rect 392 43 399 46
rect 403 43 425 46
rect 445 43 452 46
rect 466 43 471 46
rect 475 43 499 46
rect 524 43 531 46
rect 535 43 557 46
rect 218 33 225 36
rect 229 37 248 40
rect 248 30 251 36
rect 276 33 283 36
rect 287 37 302 40
rect 350 33 357 36
rect 361 37 380 40
rect 380 30 383 36
rect 408 33 415 36
rect 419 37 434 40
rect 482 33 489 36
rect 493 37 512 40
rect 512 30 515 36
rect 540 33 547 36
rect 551 37 568 40
rect 185 14 188 26
rect 206 14 209 26
rect 222 14 225 26
rect 236 17 248 20
rect 264 14 267 26
rect 280 14 283 26
rect 301 14 304 26
rect 317 14 320 26
rect 338 14 341 26
rect 354 14 357 26
rect 368 17 380 20
rect 396 14 399 26
rect 412 14 415 26
rect 433 14 436 26
rect 449 14 452 26
rect 470 14 473 26
rect 486 14 489 26
rect 500 17 512 20
rect 528 14 531 26
rect 544 14 547 26
rect 565 14 568 26
rect 182 10 215 14
rect 219 10 243 14
rect 247 10 273 14
rect 277 10 347 14
rect 351 10 375 14
rect 379 10 405 14
rect 409 10 479 14
rect 483 10 507 14
rect 511 10 537 14
rect 541 10 594 14
rect 182 3 191 7
rect 195 3 242 7
rect 246 3 292 7
rect 296 3 323 7
rect 327 3 374 7
rect 378 3 424 7
rect 428 3 455 7
rect 459 3 506 7
rect 510 3 556 7
rect 560 3 630 7
<< m2contact >>
rect 642 975 648 979
rect 663 975 667 979
rect 699 975 703 979
rect 766 975 770 979
rect 795 975 799 979
rect 831 975 835 979
rect 898 975 902 979
rect 927 975 931 979
rect 963 975 967 979
rect 1030 975 1034 979
rect 1059 975 1063 979
rect 1095 975 1099 979
rect 1162 975 1166 979
rect 582 968 588 972
rect 663 961 667 965
rect 713 961 717 965
rect 766 961 770 965
rect 795 961 799 965
rect 845 961 849 965
rect 898 961 902 965
rect 927 961 931 965
rect 977 961 981 965
rect 1030 961 1034 965
rect 1059 961 1063 965
rect 1109 961 1113 965
rect 1162 961 1166 965
rect 686 950 690 954
rect 323 942 327 946
rect 359 942 363 946
rect 426 942 430 946
rect 642 942 648 946
rect 657 941 661 945
rect 670 944 674 950
rect 707 944 711 950
rect 720 946 724 950
rect 744 950 748 954
rect 818 950 822 954
rect 728 944 732 950
rect 765 944 769 950
rect 781 946 785 950
rect 582 935 588 939
rect 323 928 327 932
rect 373 928 377 932
rect 426 928 430 932
rect 670 931 674 935
rect 686 931 690 937
rect 720 937 724 941
rect 707 931 711 935
rect 728 931 732 935
rect 744 931 748 937
rect 789 941 793 945
rect 802 944 806 950
rect 839 944 843 950
rect 852 946 856 950
rect 876 950 880 954
rect 950 950 954 954
rect 860 944 864 950
rect 897 944 901 950
rect 913 946 917 950
rect 765 931 769 935
rect 781 931 785 935
rect 802 931 806 935
rect 818 931 822 937
rect 852 937 856 941
rect 839 931 843 935
rect 860 931 864 935
rect 876 931 880 937
rect 921 941 925 945
rect 934 944 938 950
rect 971 944 975 950
rect 984 946 988 950
rect 1008 950 1012 954
rect 1082 950 1086 954
rect 992 944 996 950
rect 1029 944 1033 950
rect 1045 946 1049 950
rect 897 931 901 935
rect 913 931 917 935
rect 934 931 938 935
rect 950 931 954 937
rect 984 937 988 941
rect 971 931 975 935
rect 992 931 996 935
rect 1008 931 1012 937
rect 1053 941 1057 945
rect 1066 944 1070 950
rect 1103 944 1107 950
rect 1116 946 1120 950
rect 1140 950 1144 954
rect 1124 944 1128 950
rect 1161 944 1165 950
rect 1177 946 1181 950
rect 1029 931 1033 935
rect 1045 931 1049 935
rect 1066 931 1070 935
rect 1082 931 1086 937
rect 1116 937 1120 941
rect 1103 931 1107 935
rect 346 917 350 921
rect 308 908 312 912
rect 330 911 334 917
rect 367 911 371 917
rect 380 913 384 917
rect 404 917 408 921
rect 388 911 392 917
rect 425 911 429 917
rect 441 911 445 917
rect 663 920 667 924
rect 700 918 704 922
rect 720 918 724 922
rect 764 918 768 922
rect 795 920 799 924
rect 832 918 836 922
rect 852 918 856 922
rect 896 918 900 922
rect 927 920 931 924
rect 964 918 968 922
rect 984 918 988 922
rect 1028 918 1032 922
rect 1045 923 1049 927
rect 1124 931 1128 935
rect 1140 931 1144 937
rect 1161 931 1165 935
rect 1177 931 1181 935
rect 1059 920 1063 924
rect 1096 918 1100 922
rect 1116 918 1120 922
rect 1160 918 1164 922
rect 1177 923 1181 927
rect 594 911 600 915
rect 330 898 334 902
rect 346 898 350 904
rect 380 904 384 908
rect 367 898 371 902
rect 388 898 392 902
rect 404 898 408 904
rect 630 904 636 908
rect 663 904 667 908
rect 714 904 718 908
rect 764 904 768 908
rect 795 904 799 908
rect 846 904 850 908
rect 896 904 900 908
rect 927 904 931 908
rect 978 904 982 908
rect 1028 904 1032 908
rect 1059 904 1063 908
rect 1110 904 1114 908
rect 1160 904 1164 908
rect 425 898 429 902
rect 441 898 445 902
rect 323 887 327 891
rect 360 885 364 889
rect 380 885 384 889
rect 424 885 428 889
rect 582 891 588 895
rect 661 891 665 895
rect 695 891 699 895
rect 712 891 716 895
rect 768 891 772 895
rect 785 891 789 895
rect 813 891 817 895
rect 618 884 624 888
rect 688 884 692 888
rect 719 884 723 888
rect 741 884 745 888
rect 806 884 810 888
rect 594 878 600 882
rect 323 871 327 875
rect 374 871 378 875
rect 424 871 428 875
rect 630 871 636 875
rect 662 874 666 878
rect 687 877 691 881
rect 694 874 698 878
rect 712 874 716 878
rect 734 877 738 881
rect 759 877 763 881
rect 769 874 773 878
rect 785 874 789 878
rect 805 877 809 881
rect 812 874 816 878
rect 876 884 880 888
rect 441 864 445 868
rect 308 855 312 859
rect 433 857 437 861
rect 457 857 461 861
rect 316 848 320 852
rect 457 848 461 852
rect 689 858 693 862
rect 709 855 713 859
rect 728 859 732 863
rect 830 870 834 874
rect 845 870 849 874
rect 747 858 751 862
rect 766 858 770 862
rect 779 857 783 861
rect 801 858 805 862
rect 809 857 813 861
rect 821 857 825 861
rect 662 844 666 848
rect 694 844 698 848
rect 712 844 716 848
rect 769 844 773 848
rect 784 844 788 848
rect 812 844 816 848
rect 323 840 327 844
rect 390 840 394 844
rect 426 840 430 844
rect 642 840 648 844
rect 676 840 680 844
rect 719 839 723 843
rect 741 840 748 844
rect 791 839 795 843
rect 582 833 588 837
rect 323 826 327 830
rect 376 826 380 830
rect 426 826 430 830
rect 606 832 612 836
rect 676 832 680 836
rect 735 832 739 836
rect 760 832 764 836
rect 791 832 795 836
rect 884 862 888 870
rect 957 884 961 888
rect 911 870 915 874
rect 926 870 930 874
rect 907 862 911 866
rect 853 856 857 860
rect 866 848 870 852
rect 965 862 969 870
rect 992 862 996 866
rect 934 856 938 860
rect 947 848 951 852
rect 594 825 600 829
rect 662 825 666 829
rect 676 825 680 829
rect 694 825 698 829
rect 712 825 716 829
rect 735 825 739 829
rect 769 825 773 829
rect 784 825 788 829
rect 812 825 816 829
rect 345 815 349 819
rect 308 809 312 815
rect 324 809 328 815
rect 361 809 365 815
rect 369 811 373 815
rect 403 815 407 819
rect 606 818 612 822
rect 676 818 680 822
rect 735 818 739 822
rect 760 818 764 822
rect 791 818 795 822
rect 382 809 386 815
rect 419 809 423 815
rect 676 810 680 814
rect 719 811 723 815
rect 741 810 748 814
rect 791 811 795 815
rect 441 806 445 810
rect 662 806 666 810
rect 694 806 698 810
rect 712 806 716 810
rect 769 806 773 810
rect 784 806 788 810
rect 812 806 816 810
rect 308 796 312 800
rect 324 796 328 800
rect 369 802 373 806
rect 345 796 349 802
rect 361 796 365 800
rect 382 796 386 800
rect 403 796 407 802
rect 419 796 423 800
rect 657 794 661 798
rect 325 783 329 787
rect 369 783 373 787
rect 389 783 393 787
rect 426 785 430 789
rect 689 792 693 796
rect 709 795 713 799
rect 728 791 732 795
rect 747 792 751 796
rect 766 792 770 796
rect 779 793 783 797
rect 876 808 880 812
rect 957 808 961 812
rect 801 792 805 796
rect 809 793 813 797
rect 821 793 825 797
rect 856 793 860 797
rect 884 792 888 796
rect 936 793 940 797
rect 965 792 969 796
rect 594 776 600 780
rect 662 776 666 780
rect 687 773 691 777
rect 694 776 698 780
rect 712 776 716 780
rect 734 773 738 777
rect 759 773 763 777
rect 769 776 773 780
rect 785 776 789 780
rect 805 773 809 777
rect 812 776 816 780
rect 325 769 329 773
rect 375 769 379 773
rect 426 769 430 773
rect 630 769 636 773
rect 672 766 676 770
rect 688 766 692 770
rect 719 766 723 770
rect 741 766 745 770
rect 806 766 810 770
rect 866 772 870 776
rect 947 772 951 776
rect 582 759 588 763
rect 661 759 665 763
rect 695 759 699 763
rect 712 759 716 763
rect 768 759 772 763
rect 785 759 789 763
rect 813 759 817 763
rect 618 752 624 756
rect 672 752 676 756
rect 688 752 692 756
rect 719 752 723 756
rect 741 752 745 756
rect 806 752 810 756
rect 876 752 880 756
rect 662 742 666 746
rect 687 745 691 749
rect 694 742 698 746
rect 712 742 716 746
rect 734 745 738 749
rect 759 745 763 749
rect 769 742 773 746
rect 785 742 789 746
rect 805 745 809 749
rect 812 742 816 746
rect 656 725 660 729
rect 689 726 693 730
rect 709 723 713 727
rect 728 727 732 731
rect 747 726 751 730
rect 766 726 770 730
rect 779 725 783 729
rect 801 726 805 730
rect 809 725 813 729
rect 821 725 825 729
rect 884 730 888 738
rect 981 752 985 756
rect 935 738 939 742
rect 950 738 954 742
rect 853 724 857 728
rect 907 729 911 733
rect 662 712 666 716
rect 694 712 698 716
rect 712 712 716 716
rect 769 712 773 716
rect 784 712 788 716
rect 812 712 816 716
rect 676 708 680 712
rect 719 707 723 711
rect 741 708 748 712
rect 791 707 795 711
rect 606 700 612 704
rect 676 700 680 704
rect 735 700 739 704
rect 760 700 764 704
rect 791 700 795 704
rect 866 716 870 720
rect 989 730 993 738
rect 1010 730 1014 734
rect 958 724 962 728
rect 971 716 975 720
rect 594 693 600 697
rect 662 693 666 697
rect 676 693 680 697
rect 694 693 698 697
rect 712 693 716 697
rect 735 693 739 697
rect 769 693 773 697
rect 784 693 788 697
rect 812 693 816 697
rect 606 686 612 690
rect 676 686 680 690
rect 735 686 739 690
rect 760 686 764 690
rect 791 686 795 690
rect 676 678 680 682
rect 719 679 723 683
rect 741 678 748 682
rect 791 679 795 683
rect 662 674 666 678
rect 694 674 698 678
rect 712 674 716 678
rect 769 674 773 678
rect 784 674 788 678
rect 812 674 816 678
rect 876 677 880 681
rect 981 677 985 681
rect 657 662 661 666
rect 689 660 693 664
rect 709 663 713 667
rect 728 659 732 663
rect 747 660 751 664
rect 766 660 770 664
rect 779 661 783 665
rect 801 660 805 664
rect 809 661 813 665
rect 821 661 825 665
rect 855 662 859 666
rect 884 661 888 665
rect 961 662 965 666
rect 989 661 993 665
rect 662 644 666 648
rect 687 641 691 645
rect 694 644 698 648
rect 712 644 716 648
rect 734 641 738 645
rect 759 641 763 645
rect 769 644 773 648
rect 785 644 789 648
rect 805 641 809 645
rect 812 644 816 648
rect 618 634 624 638
rect 688 634 692 638
rect 719 634 723 638
rect 741 634 745 638
rect 806 634 810 638
rect 866 641 870 645
rect 971 641 975 645
rect 582 627 588 631
rect 661 627 665 631
rect 695 627 699 631
rect 712 627 716 631
rect 768 627 772 631
rect 785 627 789 631
rect 813 627 817 631
rect 618 620 624 624
rect 688 620 692 624
rect 719 620 723 624
rect 741 620 745 624
rect 806 620 810 624
rect 876 620 880 624
rect 662 610 666 614
rect 687 613 691 617
rect 694 610 698 614
rect 712 610 716 614
rect 734 613 738 617
rect 759 613 763 617
rect 769 610 773 614
rect 785 610 789 614
rect 805 613 809 617
rect 812 610 816 614
rect 656 593 660 597
rect 689 594 693 598
rect 709 591 713 595
rect 728 595 732 599
rect 747 594 751 598
rect 766 594 770 598
rect 779 593 783 597
rect 801 594 805 598
rect 809 593 813 597
rect 821 593 825 597
rect 884 598 888 606
rect 957 620 961 624
rect 911 606 915 610
rect 926 606 930 610
rect 907 598 911 602
rect 853 592 857 596
rect 662 580 666 584
rect 694 580 698 584
rect 712 580 716 584
rect 769 580 773 584
rect 784 580 788 584
rect 812 580 816 584
rect 676 576 680 580
rect 719 575 723 579
rect 741 576 748 580
rect 791 575 795 579
rect 606 568 612 572
rect 676 568 680 572
rect 735 568 739 572
rect 760 568 764 572
rect 791 568 795 572
rect 866 584 870 588
rect 965 598 969 606
rect 1047 620 1051 624
rect 1001 606 1005 610
rect 1016 606 1020 610
rect 989 598 993 602
rect 934 592 938 596
rect 1023 600 1027 604
rect 1055 598 1059 606
rect 947 584 951 588
rect 1090 597 1094 601
rect 1037 584 1041 588
rect 594 561 600 565
rect 662 561 666 565
rect 676 561 680 565
rect 694 561 698 565
rect 712 561 716 565
rect 735 561 739 565
rect 769 561 773 565
rect 784 561 788 565
rect 812 561 816 565
rect 606 554 612 558
rect 676 554 680 558
rect 735 554 739 558
rect 760 554 764 558
rect 791 554 795 558
rect 676 546 680 550
rect 719 547 723 551
rect 741 546 748 550
rect 791 547 795 551
rect 662 542 666 546
rect 694 542 698 546
rect 712 542 716 546
rect 769 542 773 546
rect 784 542 788 546
rect 812 542 816 546
rect 657 530 661 534
rect 689 528 693 532
rect 709 531 713 535
rect 728 527 732 531
rect 747 528 751 532
rect 766 528 770 532
rect 779 529 783 533
rect 876 542 880 546
rect 957 542 961 546
rect 1047 542 1051 546
rect 801 528 805 532
rect 809 529 813 533
rect 821 529 825 533
rect 856 527 860 531
rect 884 526 888 530
rect 936 527 940 531
rect 965 526 969 530
rect 1020 527 1024 531
rect 1055 526 1059 530
rect 662 512 666 516
rect 687 509 691 513
rect 694 512 698 516
rect 712 512 716 516
rect 734 509 738 513
rect 759 509 763 513
rect 769 512 773 516
rect 785 512 789 516
rect 805 509 809 513
rect 812 512 816 516
rect 618 502 624 506
rect 688 502 692 506
rect 719 502 723 506
rect 741 502 745 506
rect 806 502 810 506
rect 866 506 870 510
rect 947 506 951 510
rect 1037 506 1041 510
rect 582 495 588 499
rect 661 495 665 499
rect 695 495 699 499
rect 712 495 716 499
rect 768 495 772 499
rect 785 495 789 499
rect 813 495 817 499
rect 618 488 624 492
rect 688 488 692 492
rect 719 488 723 492
rect 741 488 745 492
rect 806 488 810 492
rect 876 488 880 492
rect 662 478 666 482
rect 687 481 691 485
rect 694 478 698 482
rect 712 478 716 482
rect 734 481 738 485
rect 759 481 763 485
rect 769 478 773 482
rect 785 478 789 482
rect 805 481 809 485
rect 812 478 816 482
rect 656 461 660 465
rect 689 462 693 466
rect 709 459 713 463
rect 728 463 732 467
rect 747 462 751 466
rect 766 462 770 466
rect 779 461 783 465
rect 801 462 805 466
rect 809 461 813 465
rect 821 461 825 465
rect 884 466 888 474
rect 853 460 857 464
rect 907 465 911 469
rect 662 448 666 452
rect 694 448 698 452
rect 712 448 716 452
rect 769 448 773 452
rect 784 448 788 452
rect 812 448 816 452
rect 676 444 680 448
rect 191 440 195 444
rect 227 440 231 444
rect 294 440 298 444
rect 323 440 327 444
rect 359 440 363 444
rect 426 440 430 444
rect 455 440 459 444
rect 491 440 495 444
rect 558 440 562 444
rect 642 440 648 444
rect 719 443 723 447
rect 741 444 748 448
rect 791 443 795 447
rect 582 433 588 437
rect 676 436 680 440
rect 685 436 689 440
rect 735 436 739 440
rect 760 436 764 440
rect 791 436 795 440
rect 866 452 870 456
rect 191 426 195 430
rect 241 426 245 430
rect 294 426 298 430
rect 323 426 327 430
rect 373 426 377 430
rect 426 426 430 430
rect 455 426 459 430
rect 505 426 509 430
rect 558 426 562 430
rect 594 429 600 433
rect 662 429 666 433
rect 676 429 680 433
rect 694 429 698 433
rect 712 429 716 433
rect 735 429 739 433
rect 769 429 773 433
rect 784 429 788 433
rect 812 429 816 433
rect 937 429 941 433
rect 955 429 959 433
rect 973 429 977 433
rect 996 429 1000 433
rect 1030 429 1034 433
rect 1045 429 1049 433
rect 1073 429 1077 433
rect 214 415 218 419
rect 185 406 189 410
rect 198 409 202 415
rect 235 409 239 415
rect 248 411 252 415
rect 272 415 276 419
rect 346 415 350 419
rect 256 409 260 415
rect 293 409 297 415
rect 309 409 313 415
rect 330 409 334 415
rect 367 409 371 415
rect 380 411 384 415
rect 404 415 408 419
rect 478 415 482 419
rect 388 409 392 415
rect 425 409 429 415
rect 441 409 445 415
rect 462 409 466 415
rect 499 409 503 415
rect 512 411 516 415
rect 536 415 540 419
rect 606 422 612 426
rect 676 422 680 426
rect 685 422 689 426
rect 735 422 739 426
rect 760 422 764 426
rect 791 422 795 426
rect 520 409 524 415
rect 557 409 561 415
rect 573 411 577 415
rect 676 414 680 418
rect 719 415 723 419
rect 741 414 748 418
rect 791 415 795 419
rect 662 410 666 414
rect 694 410 698 414
rect 712 410 716 414
rect 769 410 773 414
rect 784 410 788 414
rect 812 410 816 414
rect 198 396 202 400
rect 214 396 218 402
rect 248 402 252 406
rect 235 396 239 400
rect 256 396 260 400
rect 272 396 276 402
rect 293 396 297 400
rect 309 396 313 400
rect 330 396 334 400
rect 346 396 350 402
rect 380 402 384 406
rect 367 396 371 400
rect 388 396 392 400
rect 404 396 408 402
rect 425 396 429 400
rect 441 396 445 400
rect 462 396 466 400
rect 478 396 482 402
rect 512 402 516 406
rect 499 396 503 400
rect 520 396 524 400
rect 536 396 540 402
rect 557 396 561 400
rect 573 396 577 400
rect 657 398 661 402
rect 191 385 195 389
rect 228 383 232 387
rect 248 383 252 387
rect 292 383 296 387
rect 323 385 327 389
rect 360 383 364 387
rect 380 383 384 387
rect 424 383 428 387
rect 455 385 459 389
rect 492 383 496 387
rect 512 383 516 387
rect 556 383 560 387
rect 689 396 693 400
rect 709 399 713 403
rect 728 395 732 399
rect 747 396 751 400
rect 766 396 770 400
rect 779 397 783 401
rect 915 422 919 426
rect 937 422 941 426
rect 996 422 1000 426
rect 1021 422 1025 426
rect 1052 422 1056 426
rect 937 414 941 418
rect 980 415 984 419
rect 1002 414 1009 418
rect 1052 415 1056 419
rect 955 410 959 414
rect 973 410 977 414
rect 1030 410 1034 414
rect 1045 410 1049 414
rect 1073 410 1077 414
rect 876 406 880 410
rect 801 396 805 400
rect 809 397 813 401
rect 821 397 825 401
rect 855 391 859 395
rect 895 397 899 401
rect 884 390 888 394
rect 662 380 666 384
rect 594 376 600 380
rect 687 377 691 381
rect 694 380 698 384
rect 712 380 716 384
rect 734 377 738 381
rect 759 377 763 381
rect 769 380 773 384
rect 785 380 789 384
rect 805 377 809 381
rect 812 380 816 384
rect 950 396 954 400
rect 970 399 974 403
rect 989 395 993 399
rect 1008 396 1012 400
rect 1027 396 1031 400
rect 1040 397 1044 401
rect 1062 396 1066 400
rect 1070 397 1074 401
rect 1082 397 1086 401
rect 896 380 900 384
rect 922 380 926 384
rect 191 369 195 373
rect 242 369 246 373
rect 292 369 296 373
rect 323 369 327 373
rect 374 369 378 373
rect 424 369 428 373
rect 455 369 459 373
rect 506 369 510 373
rect 556 369 560 373
rect 630 370 636 374
rect 670 370 674 374
rect 688 370 692 374
rect 719 370 723 374
rect 741 370 745 374
rect 806 370 810 374
rect 948 377 952 381
rect 955 380 959 384
rect 973 380 977 384
rect 995 377 999 381
rect 1020 377 1024 381
rect 1030 380 1034 384
rect 1046 380 1050 384
rect 1066 377 1070 381
rect 1073 380 1077 384
rect 866 370 870 374
rect 905 370 909 374
rect 949 370 953 374
rect 980 370 984 374
rect 1002 370 1006 374
rect 1067 370 1071 374
rect 185 362 189 366
rect 573 362 577 366
rect 582 363 588 367
rect 661 363 665 367
rect 695 363 699 367
rect 712 363 716 367
rect 768 363 772 367
rect 785 363 789 367
rect 813 363 817 367
rect 896 363 900 367
rect 922 363 926 367
rect 956 363 960 367
rect 973 363 977 367
rect 1029 363 1033 367
rect 1046 363 1050 367
rect 1074 363 1078 367
rect 308 355 313 359
rect 441 355 445 359
rect 618 356 624 360
rect 670 356 674 360
rect 904 356 908 360
rect 1090 357 1094 361
rect 1102 357 1106 361
rect 316 348 320 352
rect 606 348 612 352
rect 914 349 918 353
rect 1079 349 1083 353
rect 300 344 304 348
rect 332 344 336 348
rect 300 337 304 341
rect 332 337 336 341
rect 316 330 320 334
rect 573 330 577 334
rect 642 330 648 334
rect 962 330 966 334
rect 998 330 1002 334
rect 1065 330 1069 334
rect 573 322 577 326
rect 582 323 588 327
rect 948 323 952 327
rect 300 318 304 322
rect 332 318 336 322
rect 316 314 320 318
rect 962 316 966 320
rect 1012 316 1016 320
rect 1065 316 1069 320
rect 308 307 313 311
rect 442 307 446 311
rect 985 305 989 309
rect 191 300 195 304
rect 227 300 231 304
rect 294 300 298 304
rect 323 300 327 304
rect 359 300 363 304
rect 426 300 430 304
rect 455 300 459 304
rect 491 300 495 304
rect 558 300 562 304
rect 642 300 648 304
rect 582 293 588 297
rect 956 296 960 300
rect 969 299 973 305
rect 1006 299 1010 305
rect 1019 301 1023 305
rect 1043 305 1047 309
rect 1027 299 1031 305
rect 1064 299 1068 305
rect 1080 299 1084 305
rect 191 286 195 290
rect 241 286 245 290
rect 294 286 298 290
rect 323 286 327 290
rect 373 286 377 290
rect 426 286 430 290
rect 455 286 459 290
rect 505 286 509 290
rect 558 286 562 290
rect 969 286 973 290
rect 985 286 989 292
rect 1019 292 1023 296
rect 1006 286 1010 290
rect 214 275 218 279
rect 185 266 189 270
rect 198 269 202 275
rect 235 269 239 275
rect 248 271 252 275
rect 272 275 276 279
rect 346 275 350 279
rect 256 269 260 275
rect 293 269 297 275
rect 309 269 313 275
rect 330 269 334 275
rect 367 269 371 275
rect 380 271 384 275
rect 404 275 408 279
rect 478 275 482 279
rect 388 269 392 275
rect 425 269 429 275
rect 441 269 445 275
rect 462 269 466 275
rect 499 269 503 275
rect 512 271 516 275
rect 536 275 540 279
rect 520 269 524 275
rect 557 269 561 275
rect 573 271 577 275
rect 1027 286 1031 290
rect 1043 286 1047 292
rect 1064 286 1068 290
rect 1080 286 1084 290
rect 962 275 966 279
rect 999 273 1003 277
rect 1019 273 1023 277
rect 1063 273 1067 277
rect 198 256 202 260
rect 214 256 218 262
rect 248 262 252 266
rect 235 256 239 260
rect 256 256 260 260
rect 272 256 276 262
rect 293 256 297 260
rect 309 256 313 260
rect 330 256 334 260
rect 346 256 350 262
rect 380 262 384 266
rect 367 256 371 260
rect 388 256 392 260
rect 404 256 408 262
rect 425 256 429 260
rect 441 256 445 260
rect 462 256 466 260
rect 478 256 482 262
rect 512 262 516 266
rect 499 256 503 260
rect 520 256 524 260
rect 536 256 540 262
rect 594 266 600 270
rect 557 256 561 260
rect 573 256 577 260
rect 630 259 636 263
rect 962 259 966 263
rect 1013 259 1017 263
rect 1063 259 1067 263
rect 191 245 195 249
rect 228 243 232 247
rect 248 243 252 247
rect 292 243 296 247
rect 323 245 327 249
rect 360 243 364 247
rect 380 243 384 247
rect 424 243 428 247
rect 455 245 459 249
rect 492 243 496 247
rect 512 243 516 247
rect 556 243 560 247
rect 955 251 959 255
rect 1080 252 1084 256
rect 642 244 648 248
rect 962 244 966 248
rect 998 244 1002 248
rect 1065 244 1069 248
rect 594 236 600 240
rect 948 237 952 241
rect 191 229 195 233
rect 242 229 246 233
rect 292 229 296 233
rect 323 229 327 233
rect 374 229 378 233
rect 424 229 428 233
rect 455 229 459 233
rect 506 229 510 233
rect 556 229 560 233
rect 630 229 636 233
rect 962 230 966 234
rect 1012 230 1016 234
rect 1065 230 1069 234
rect 184 222 188 226
rect 573 222 577 226
rect 985 219 989 223
rect 191 214 195 218
rect 227 214 231 218
rect 294 214 298 218
rect 323 214 327 218
rect 359 214 363 218
rect 426 214 430 218
rect 455 214 459 218
rect 491 214 495 218
rect 558 214 562 218
rect 642 214 648 218
rect 582 207 588 211
rect 956 210 960 214
rect 969 213 973 219
rect 1006 213 1010 219
rect 1019 215 1023 219
rect 1043 219 1047 223
rect 1027 213 1031 219
rect 1064 213 1068 219
rect 1080 215 1084 219
rect 1102 213 1106 217
rect 191 200 195 204
rect 241 200 245 204
rect 294 200 298 204
rect 323 200 327 204
rect 373 200 377 204
rect 426 200 430 204
rect 455 200 459 204
rect 505 200 509 204
rect 558 200 562 204
rect 969 200 973 204
rect 985 200 989 206
rect 1019 206 1023 210
rect 1006 200 1010 204
rect 214 189 218 193
rect 185 180 189 184
rect 198 183 202 189
rect 235 183 239 189
rect 248 185 252 189
rect 272 189 276 193
rect 346 189 350 193
rect 256 183 260 189
rect 293 183 297 189
rect 309 183 313 189
rect 330 183 334 189
rect 367 183 371 189
rect 380 185 384 189
rect 404 189 408 193
rect 478 189 482 193
rect 388 183 392 189
rect 425 183 429 189
rect 441 183 445 189
rect 462 183 466 189
rect 499 183 503 189
rect 512 185 516 189
rect 536 189 540 193
rect 520 183 524 189
rect 557 183 561 189
rect 573 185 577 189
rect 1027 200 1031 204
rect 1043 200 1047 206
rect 1064 200 1068 204
rect 1080 200 1084 209
rect 1102 197 1106 201
rect 962 189 966 193
rect 999 187 1003 191
rect 1019 187 1023 191
rect 1063 187 1067 191
rect 198 170 202 174
rect 214 170 218 176
rect 248 176 252 180
rect 235 170 239 174
rect 256 170 260 174
rect 272 170 276 176
rect 293 170 297 174
rect 309 170 313 174
rect 330 170 334 174
rect 346 170 350 176
rect 380 176 384 180
rect 367 170 371 174
rect 388 170 392 174
rect 404 170 408 176
rect 425 170 429 174
rect 441 170 445 174
rect 462 170 466 174
rect 478 170 482 176
rect 512 176 516 180
rect 499 170 503 174
rect 520 170 524 174
rect 536 170 540 176
rect 594 180 600 184
rect 557 170 561 174
rect 573 170 577 174
rect 630 173 636 177
rect 962 173 966 177
rect 1013 173 1017 177
rect 1063 173 1067 177
rect 191 159 195 163
rect 228 157 232 161
rect 248 157 252 161
rect 292 157 296 161
rect 323 159 327 163
rect 360 157 364 161
rect 380 157 384 161
rect 424 157 428 161
rect 455 159 459 163
rect 492 157 496 161
rect 512 157 516 161
rect 556 157 560 161
rect 594 150 600 154
rect 191 143 195 147
rect 242 143 246 147
rect 292 143 296 147
rect 323 143 327 147
rect 374 143 378 147
rect 424 143 428 147
rect 455 143 459 147
rect 506 143 510 147
rect 556 143 560 147
rect 630 143 636 147
rect 184 136 188 140
rect 573 136 577 140
rect 309 129 313 133
rect 417 129 421 133
rect 441 129 445 133
rect 433 122 437 126
rect 417 118 421 122
rect 449 118 453 122
rect 417 111 421 115
rect 449 111 453 115
rect 1102 111 1106 115
rect 433 104 437 108
rect 573 104 577 108
rect 573 96 577 100
rect 417 92 421 96
rect 449 92 453 96
rect 433 88 437 92
rect 309 81 313 85
rect 417 81 421 85
rect 441 81 445 85
rect 191 74 195 78
rect 227 74 231 78
rect 294 74 298 78
rect 323 74 327 78
rect 359 74 363 78
rect 426 74 430 78
rect 455 74 459 78
rect 491 74 495 78
rect 558 74 562 78
rect 642 74 648 78
rect 582 67 588 71
rect 191 60 195 64
rect 241 60 245 64
rect 294 60 298 64
rect 323 60 327 64
rect 373 60 377 64
rect 426 60 430 64
rect 455 60 459 64
rect 505 60 509 64
rect 558 60 562 64
rect 214 49 218 53
rect 185 40 189 44
rect 198 43 202 49
rect 235 43 239 49
rect 248 45 252 49
rect 272 49 276 53
rect 346 49 350 53
rect 256 43 260 49
rect 293 43 297 49
rect 309 43 313 49
rect 330 43 334 49
rect 367 43 371 49
rect 380 45 384 49
rect 404 49 408 53
rect 478 49 482 53
rect 388 43 392 49
rect 425 43 429 49
rect 441 43 445 49
rect 462 43 466 49
rect 499 43 503 49
rect 512 45 516 49
rect 536 49 540 53
rect 520 43 524 49
rect 557 43 561 49
rect 573 45 577 49
rect 198 30 202 34
rect 214 30 218 36
rect 248 36 252 40
rect 235 30 239 34
rect 256 30 260 34
rect 272 30 276 36
rect 293 30 297 34
rect 309 30 313 34
rect 330 30 334 34
rect 346 30 350 36
rect 380 36 384 40
rect 367 30 371 34
rect 388 30 392 34
rect 404 30 408 36
rect 425 30 429 34
rect 441 30 445 34
rect 462 30 466 34
rect 478 30 482 36
rect 512 36 516 40
rect 499 30 503 34
rect 520 30 524 34
rect 536 30 540 36
rect 557 30 561 34
rect 573 30 577 34
rect 191 19 195 23
rect 228 17 232 21
rect 248 17 252 21
rect 292 17 296 21
rect 323 19 327 23
rect 360 17 364 21
rect 380 17 384 21
rect 424 17 428 21
rect 455 19 459 23
rect 492 17 496 21
rect 512 17 516 21
rect 556 17 560 21
rect 594 10 600 14
rect 191 3 195 7
rect 242 3 246 7
rect 292 3 296 7
rect 323 3 327 7
rect 374 3 378 7
rect 424 3 428 7
rect 455 3 459 7
rect 506 3 510 7
rect 556 3 560 7
rect 630 3 636 7
<< metal2 >>
rect 308 859 311 908
rect 308 815 311 855
rect 316 852 320 995
rect 324 932 327 942
rect 331 902 334 911
rect 347 904 350 917
rect 360 889 363 942
rect 427 932 430 942
rect 367 917 371 921
rect 368 902 371 911
rect 323 875 326 887
rect 364 885 365 889
rect 374 875 377 928
rect 380 908 383 913
rect 389 902 392 911
rect 405 904 408 917
rect 426 902 429 911
rect 425 875 428 885
rect 308 800 311 809
rect 192 430 195 440
rect 199 400 202 409
rect 215 402 218 415
rect 228 387 231 440
rect 295 430 298 440
rect 235 415 239 419
rect 236 400 239 409
rect 191 373 194 385
rect 232 383 233 387
rect 242 373 245 426
rect 248 406 251 411
rect 257 400 260 409
rect 273 402 276 415
rect 294 400 297 409
rect 310 400 313 409
rect 293 373 296 383
rect 185 270 188 362
rect 310 359 313 396
rect 316 352 320 848
rect 433 861 437 995
rect 582 972 588 986
rect 582 939 588 968
rect 442 909 445 911
rect 442 902 445 905
rect 442 868 445 898
rect 582 895 588 935
rect 323 830 326 840
rect 324 800 327 809
rect 345 802 348 815
rect 361 800 364 809
rect 370 806 373 811
rect 325 773 328 783
rect 376 773 379 826
rect 382 815 386 819
rect 382 800 385 809
rect 390 787 393 840
rect 426 830 429 840
rect 403 802 406 815
rect 419 800 422 809
rect 388 783 389 787
rect 427 773 430 785
rect 324 430 327 440
rect 331 400 334 409
rect 347 402 350 415
rect 360 387 363 440
rect 427 430 430 440
rect 367 415 371 419
rect 368 400 371 409
rect 323 373 326 385
rect 364 383 365 387
rect 374 373 377 426
rect 380 406 383 411
rect 389 400 392 409
rect 405 402 408 415
rect 426 400 429 409
rect 425 373 428 383
rect 300 341 304 344
rect 300 322 304 337
rect 316 334 320 348
rect 332 348 336 352
rect 332 341 336 344
rect 332 322 336 337
rect 316 318 320 319
rect 332 314 336 318
rect 192 290 195 300
rect 199 260 202 269
rect 215 262 218 275
rect 228 247 231 300
rect 295 290 298 300
rect 235 275 239 279
rect 236 260 239 269
rect 191 233 194 245
rect 232 243 233 247
rect 242 233 245 286
rect 310 275 313 307
rect 248 266 251 271
rect 257 260 260 269
rect 273 262 276 275
rect 294 260 297 269
rect 310 260 313 269
rect 293 233 296 243
rect 185 184 188 222
rect 192 204 195 214
rect 199 174 202 183
rect 215 176 218 189
rect 228 161 231 214
rect 295 204 298 214
rect 235 189 239 193
rect 236 174 239 183
rect 191 147 194 159
rect 232 157 233 161
rect 242 147 245 200
rect 248 180 251 185
rect 257 174 260 183
rect 273 176 276 189
rect 294 174 297 183
rect 310 174 313 183
rect 293 147 296 157
rect 185 44 188 136
rect 310 133 313 170
rect 192 64 195 74
rect 199 34 202 43
rect 215 36 218 49
rect 228 21 231 74
rect 295 64 298 74
rect 235 49 239 53
rect 236 34 239 43
rect 191 7 194 19
rect 232 17 233 21
rect 242 7 245 60
rect 310 49 313 81
rect 248 40 251 45
rect 257 34 260 43
rect 273 36 276 49
rect 294 34 297 43
rect 310 34 313 43
rect 293 7 296 17
rect 316 0 320 314
rect 324 290 327 300
rect 331 260 334 269
rect 347 262 350 275
rect 360 247 363 300
rect 427 290 430 300
rect 367 275 371 279
rect 368 260 371 269
rect 323 233 326 245
rect 364 243 365 247
rect 374 233 377 286
rect 380 266 383 271
rect 389 260 392 269
rect 405 262 408 275
rect 426 260 429 269
rect 425 233 428 243
rect 324 204 327 214
rect 331 174 334 183
rect 347 176 350 189
rect 360 161 363 214
rect 427 204 430 214
rect 367 189 371 193
rect 368 174 371 183
rect 323 147 326 159
rect 364 157 365 161
rect 374 147 377 200
rect 380 180 383 185
rect 389 174 392 183
rect 405 176 408 189
rect 426 174 429 183
rect 425 147 428 157
rect 433 126 437 857
rect 457 852 461 857
rect 582 837 588 891
rect 582 763 588 833
rect 582 631 588 759
rect 582 499 588 627
rect 456 430 459 440
rect 442 400 445 409
rect 463 400 466 409
rect 479 402 482 415
rect 442 359 445 396
rect 492 387 495 440
rect 559 430 562 440
rect 582 437 588 495
rect 499 415 503 419
rect 500 400 503 409
rect 455 373 458 385
rect 496 383 497 387
rect 506 373 509 426
rect 512 406 515 411
rect 521 400 524 409
rect 537 402 540 415
rect 558 400 561 409
rect 574 400 577 411
rect 557 373 560 383
rect 574 366 577 396
rect 574 334 577 362
rect 582 367 588 433
rect 582 327 588 363
rect 442 275 445 307
rect 456 290 459 300
rect 442 260 445 269
rect 463 260 466 269
rect 479 262 482 275
rect 492 247 495 300
rect 559 290 562 300
rect 499 275 503 279
rect 500 260 503 269
rect 455 233 458 245
rect 496 243 497 247
rect 506 233 509 286
rect 574 275 577 322
rect 512 266 515 271
rect 521 260 524 269
rect 537 262 540 275
rect 558 260 561 269
rect 574 260 577 271
rect 557 233 560 243
rect 574 226 577 256
rect 582 297 588 323
rect 456 204 459 214
rect 442 174 445 183
rect 463 174 466 183
rect 479 176 482 189
rect 442 133 445 170
rect 492 161 495 214
rect 559 204 562 214
rect 582 211 588 293
rect 499 189 503 193
rect 500 174 503 183
rect 455 147 458 159
rect 496 157 497 161
rect 506 147 509 200
rect 512 180 515 185
rect 521 174 524 183
rect 537 176 540 189
rect 558 174 561 183
rect 574 174 577 185
rect 557 147 560 157
rect 574 140 577 170
rect 417 115 421 118
rect 417 96 421 111
rect 433 108 437 122
rect 449 122 453 126
rect 449 115 453 118
rect 449 96 453 111
rect 574 108 577 136
rect 433 92 437 93
rect 449 88 453 92
rect 324 64 327 74
rect 331 34 334 43
rect 347 36 350 49
rect 360 21 363 74
rect 427 64 430 74
rect 367 49 371 53
rect 368 34 371 43
rect 323 7 326 19
rect 364 17 365 21
rect 374 7 377 60
rect 380 40 383 45
rect 389 34 392 43
rect 405 36 408 49
rect 426 34 429 43
rect 425 7 428 17
rect 433 0 437 88
rect 442 49 445 81
rect 456 64 459 74
rect 442 34 445 43
rect 463 34 466 43
rect 479 36 482 49
rect 492 21 495 74
rect 559 64 562 74
rect 499 49 503 53
rect 500 34 503 43
rect 455 7 458 19
rect 496 17 497 21
rect 506 7 509 60
rect 574 49 577 96
rect 512 40 515 45
rect 521 34 524 43
rect 537 36 540 49
rect 558 34 561 43
rect 574 41 577 45
rect 582 71 588 207
rect 574 34 577 37
rect 557 7 560 17
rect 582 0 588 67
rect 594 915 600 986
rect 594 882 600 911
rect 594 829 600 878
rect 594 780 600 825
rect 594 697 600 776
rect 594 565 600 693
rect 594 433 600 561
rect 594 380 600 429
rect 594 270 600 376
rect 594 240 600 266
rect 594 184 600 236
rect 594 154 600 180
rect 594 14 600 150
rect 594 0 600 10
rect 606 836 612 986
rect 606 822 612 832
rect 606 704 612 818
rect 606 690 612 700
rect 606 572 612 686
rect 606 558 612 568
rect 606 426 612 554
rect 606 352 612 422
rect 606 0 612 348
rect 618 888 624 986
rect 618 756 624 884
rect 618 638 624 752
rect 618 624 624 634
rect 618 506 624 620
rect 618 492 624 502
rect 618 360 624 488
rect 618 0 624 356
rect 630 908 636 986
rect 630 875 636 904
rect 630 773 636 871
rect 630 374 636 769
rect 630 263 636 370
rect 630 233 636 259
rect 630 177 636 229
rect 630 147 636 173
rect 630 7 636 143
rect 630 0 636 3
rect 642 979 648 986
rect 642 946 648 975
rect 664 965 667 975
rect 642 844 648 942
rect 671 935 674 944
rect 687 937 690 950
rect 700 922 703 975
rect 767 965 770 975
rect 796 965 799 975
rect 707 950 711 954
rect 708 935 711 944
rect 663 908 666 920
rect 704 918 705 922
rect 714 908 717 961
rect 720 941 723 946
rect 729 935 732 944
rect 745 937 748 950
rect 766 935 769 944
rect 782 944 785 946
rect 782 941 789 944
rect 782 935 785 941
rect 803 935 806 944
rect 819 937 822 950
rect 765 908 768 918
rect 782 901 785 931
rect 832 922 835 975
rect 899 965 902 975
rect 928 965 931 975
rect 839 950 843 954
rect 840 935 843 944
rect 795 908 798 920
rect 836 918 837 922
rect 846 908 849 961
rect 852 941 855 946
rect 861 935 864 944
rect 877 937 880 950
rect 898 935 901 944
rect 914 944 917 946
rect 914 941 921 944
rect 914 935 917 941
rect 935 935 938 944
rect 951 937 954 950
rect 897 908 900 918
rect 782 898 834 901
rect 662 878 665 891
rect 688 881 691 884
rect 695 878 698 891
rect 712 878 715 891
rect 642 444 648 840
rect 662 829 665 844
rect 676 836 679 840
rect 694 829 697 844
rect 713 829 716 844
rect 719 843 722 884
rect 735 836 738 877
rect 741 844 744 884
rect 760 836 763 877
rect 769 878 772 891
rect 785 878 788 891
rect 806 881 809 884
rect 813 878 816 891
rect 831 887 834 898
rect 914 895 917 931
rect 964 922 967 975
rect 1031 965 1034 975
rect 1060 965 1063 975
rect 971 950 975 954
rect 972 935 975 944
rect 927 908 930 920
rect 968 918 969 922
rect 978 908 981 961
rect 984 941 987 946
rect 993 935 996 944
rect 1009 937 1012 950
rect 1030 935 1033 944
rect 1046 944 1049 946
rect 1046 941 1053 944
rect 1046 935 1049 941
rect 1067 935 1070 944
rect 1083 937 1086 950
rect 1029 908 1032 918
rect 1046 901 1049 923
rect 1096 922 1099 975
rect 1163 965 1166 975
rect 1103 950 1107 954
rect 1104 935 1107 944
rect 1059 908 1062 920
rect 1100 918 1101 922
rect 1110 908 1113 961
rect 1116 941 1119 946
rect 1125 935 1128 944
rect 1141 937 1144 950
rect 1162 935 1165 944
rect 1178 944 1181 946
rect 1178 941 1182 944
rect 1178 935 1181 941
rect 1178 927 1181 931
rect 1161 908 1164 918
rect 912 890 917 895
rect 974 897 1049 901
rect 831 884 876 887
rect 831 874 834 884
rect 849 871 869 874
rect 866 852 869 871
rect 769 829 772 844
rect 784 829 787 844
rect 791 836 795 839
rect 812 829 815 844
rect 662 810 665 825
rect 676 814 679 818
rect 694 810 697 825
rect 713 810 716 825
rect 662 763 665 776
rect 688 770 691 773
rect 662 746 665 759
rect 672 756 676 766
rect 695 763 698 776
rect 712 763 715 776
rect 719 770 722 811
rect 735 777 738 818
rect 741 770 744 810
rect 760 777 763 818
rect 769 810 772 825
rect 784 810 787 825
rect 791 815 795 818
rect 812 810 815 825
rect 769 763 772 776
rect 688 749 691 752
rect 695 746 698 759
rect 712 746 715 759
rect 662 697 665 712
rect 676 704 679 708
rect 694 697 697 712
rect 713 697 716 712
rect 719 711 722 752
rect 735 704 738 745
rect 741 712 744 752
rect 760 704 763 745
rect 769 746 772 759
rect 785 763 788 776
rect 806 770 809 773
rect 813 763 816 776
rect 866 776 869 848
rect 877 812 880 884
rect 912 887 915 890
rect 912 884 957 887
rect 912 874 915 884
rect 785 746 788 759
rect 806 749 809 752
rect 813 746 816 759
rect 866 742 869 772
rect 877 756 880 808
rect 884 796 888 862
rect 872 752 876 755
rect 865 739 869 742
rect 866 720 869 739
rect 769 697 772 712
rect 784 697 787 712
rect 791 704 795 707
rect 812 697 815 712
rect 662 678 665 693
rect 676 682 679 686
rect 694 678 697 693
rect 713 678 716 693
rect 662 631 665 644
rect 688 638 691 641
rect 662 614 665 627
rect 695 631 698 644
rect 712 631 715 644
rect 719 638 722 679
rect 735 645 738 686
rect 741 638 744 678
rect 760 645 763 686
rect 769 678 772 693
rect 784 678 787 693
rect 791 683 795 686
rect 812 678 815 693
rect 769 631 772 644
rect 688 617 691 620
rect 695 614 698 627
rect 712 614 715 627
rect 662 565 665 580
rect 676 572 679 576
rect 694 565 697 580
rect 713 565 716 580
rect 719 579 722 620
rect 735 572 738 613
rect 741 580 744 620
rect 760 572 763 613
rect 769 614 772 627
rect 785 631 788 644
rect 806 638 809 641
rect 813 631 816 644
rect 866 645 869 716
rect 877 681 880 752
rect 785 614 788 627
rect 806 617 809 620
rect 813 614 816 627
rect 866 588 869 641
rect 877 624 880 677
rect 884 665 888 730
rect 872 620 876 623
rect 915 623 918 874
rect 930 871 950 874
rect 947 852 950 871
rect 947 776 950 848
rect 958 812 961 884
rect 965 796 969 862
rect 974 763 977 897
rect 1178 894 1181 923
rect 1002 891 1109 894
rect 936 759 977 763
rect 936 755 939 759
rect 936 752 981 755
rect 936 742 939 752
rect 954 739 974 742
rect 936 737 939 738
rect 971 720 974 739
rect 971 645 974 716
rect 982 681 985 752
rect 989 665 993 730
rect 769 565 772 580
rect 784 565 787 580
rect 791 572 795 575
rect 812 565 815 580
rect 662 546 665 561
rect 676 550 679 554
rect 694 546 697 561
rect 713 546 716 561
rect 662 499 665 512
rect 688 506 691 509
rect 662 482 665 495
rect 695 499 698 512
rect 712 499 715 512
rect 719 506 722 547
rect 735 513 738 554
rect 741 506 744 546
rect 760 513 763 554
rect 769 546 772 561
rect 784 546 787 561
rect 791 551 795 554
rect 812 546 815 561
rect 769 499 772 512
rect 688 485 691 488
rect 695 482 698 495
rect 712 482 715 495
rect 642 334 648 440
rect 662 433 665 448
rect 676 440 679 444
rect 662 414 665 429
rect 685 426 689 436
rect 694 433 697 448
rect 713 433 716 448
rect 719 447 722 488
rect 735 440 738 481
rect 741 448 744 488
rect 760 440 763 481
rect 769 482 772 495
rect 785 499 788 512
rect 806 506 809 509
rect 813 499 816 512
rect 866 510 869 584
rect 877 546 880 620
rect 912 620 957 623
rect 912 610 915 620
rect 930 607 950 610
rect 785 482 788 495
rect 806 485 809 488
rect 813 482 816 495
rect 866 456 869 506
rect 877 492 880 542
rect 884 530 888 598
rect 947 588 950 607
rect 947 510 950 584
rect 958 546 961 620
rect 1002 623 1005 891
rect 1113 891 1181 894
rect 1002 620 1047 623
rect 1002 610 1005 620
rect 1020 607 1040 610
rect 965 530 969 598
rect 1037 588 1040 607
rect 1037 510 1040 584
rect 1048 546 1051 620
rect 1055 530 1059 598
rect 872 488 876 491
rect 769 433 772 448
rect 784 433 787 448
rect 791 440 795 443
rect 812 433 815 448
rect 676 418 679 422
rect 694 414 697 429
rect 713 414 716 429
rect 662 367 665 380
rect 688 374 691 377
rect 670 360 674 370
rect 695 367 698 380
rect 712 367 715 380
rect 719 374 722 415
rect 735 381 738 422
rect 741 374 744 414
rect 760 381 763 422
rect 769 414 772 429
rect 784 414 787 429
rect 791 419 795 422
rect 812 414 815 429
rect 769 367 772 380
rect 785 367 788 380
rect 806 374 809 377
rect 813 367 816 380
rect 866 374 869 452
rect 877 410 880 488
rect 884 394 888 466
rect 896 367 900 380
rect 905 360 908 370
rect 915 353 918 422
rect 937 418 940 422
rect 955 414 958 429
rect 974 414 977 429
rect 922 367 926 380
rect 949 374 952 377
rect 956 367 959 380
rect 973 367 976 380
rect 980 374 983 415
rect 996 381 999 422
rect 1002 374 1005 414
rect 1021 381 1024 422
rect 1030 414 1033 429
rect 1045 414 1048 429
rect 1052 419 1056 422
rect 1073 414 1076 429
rect 1030 367 1033 380
rect 1046 367 1049 380
rect 1067 374 1070 377
rect 1074 367 1077 380
rect 1090 361 1094 597
rect 1083 349 1084 352
rect 642 304 648 330
rect 642 248 648 300
rect 642 218 648 244
rect 948 241 952 323
rect 963 320 966 330
rect 970 290 973 299
rect 986 292 989 305
rect 999 277 1002 330
rect 1066 320 1069 330
rect 1006 305 1010 309
rect 1007 290 1010 299
rect 962 263 965 275
rect 1003 273 1004 277
rect 1013 263 1016 316
rect 1081 305 1084 349
rect 1019 296 1022 301
rect 1028 290 1031 299
rect 1044 292 1047 305
rect 1065 290 1068 299
rect 1081 290 1084 299
rect 1064 263 1067 273
rect 1081 256 1084 286
rect 642 78 648 214
rect 956 214 959 251
rect 963 234 966 244
rect 970 204 973 213
rect 986 206 989 219
rect 999 191 1002 244
rect 1066 234 1069 244
rect 1006 219 1010 223
rect 1007 204 1010 213
rect 962 177 965 189
rect 1003 187 1004 191
rect 1013 177 1016 230
rect 1019 210 1022 215
rect 1028 204 1031 213
rect 1044 206 1047 219
rect 1065 204 1068 213
rect 1081 214 1084 215
rect 1102 217 1106 357
rect 1081 209 1084 210
rect 1064 177 1067 187
rect 1102 115 1106 197
rect 642 0 648 74
<< m3contact >>
rect 185 402 189 406
rect 442 905 446 909
rect 441 802 445 806
rect 574 37 578 41
rect 653 941 657 945
rect 693 858 698 863
rect 704 854 709 859
rect 727 863 732 868
rect 751 858 756 863
rect 766 862 771 868
rect 796 858 801 863
rect 825 857 830 862
rect 780 852 785 857
rect 809 852 813 857
rect 851 851 856 856
rect 657 798 662 803
rect 693 791 698 796
rect 704 795 709 800
rect 727 786 732 791
rect 751 791 756 796
rect 780 797 785 802
rect 809 797 813 802
rect 766 786 771 792
rect 796 791 801 796
rect 825 792 830 797
rect 851 792 856 797
rect 656 729 661 734
rect 693 726 698 731
rect 704 722 709 727
rect 727 731 732 736
rect 751 726 756 731
rect 907 857 912 862
rect 766 730 771 736
rect 796 726 801 731
rect 825 725 830 730
rect 780 720 785 725
rect 809 720 813 725
rect 851 719 856 724
rect 657 666 662 671
rect 693 659 698 664
rect 704 663 709 668
rect 727 654 732 659
rect 751 659 756 664
rect 780 665 785 670
rect 809 665 813 670
rect 766 654 771 660
rect 796 659 801 664
rect 825 660 830 665
rect 850 661 855 666
rect 656 597 661 602
rect 693 594 698 599
rect 704 590 709 595
rect 727 599 732 604
rect 751 594 756 599
rect 766 598 771 604
rect 796 594 801 599
rect 825 593 830 598
rect 780 588 785 593
rect 809 588 813 593
rect 851 587 856 592
rect 907 733 912 738
rect 932 851 937 856
rect 931 792 936 797
rect 992 857 997 862
rect 956 719 961 724
rect 956 661 961 666
rect 657 534 662 539
rect 693 527 698 532
rect 704 531 709 536
rect 727 522 732 527
rect 751 527 756 532
rect 780 533 785 538
rect 809 533 813 538
rect 766 522 771 528
rect 796 527 801 532
rect 825 528 830 533
rect 851 526 856 531
rect 656 465 661 470
rect 693 462 698 467
rect 704 458 709 463
rect 727 467 732 472
rect 751 462 756 467
rect 766 466 771 472
rect 796 462 801 467
rect 825 461 830 466
rect 780 456 785 461
rect 809 456 813 461
rect 851 455 856 460
rect 907 593 912 598
rect 932 587 937 592
rect 931 526 936 531
rect 1109 890 1113 894
rect 1014 730 1019 735
rect 989 602 994 607
rect 1023 595 1028 600
rect 1020 522 1025 527
rect 657 402 662 407
rect 693 395 698 400
rect 704 399 709 404
rect 727 390 732 395
rect 751 395 756 400
rect 780 401 785 406
rect 809 401 813 406
rect 766 390 771 396
rect 796 395 801 400
rect 825 396 830 401
rect 850 390 855 395
rect 907 469 912 474
rect 895 401 900 406
rect 954 395 959 400
rect 965 399 970 404
rect 988 390 993 395
rect 1012 395 1017 400
rect 1041 401 1046 406
rect 1070 401 1074 406
rect 1027 390 1032 396
rect 1057 395 1062 400
rect 1082 401 1087 406
rect 956 292 960 296
rect 1081 210 1085 214
<< metal3 >>
rect 652 945 658 946
rect 652 941 653 945
rect 657 941 658 945
rect 652 940 658 941
rect 652 910 657 940
rect 441 909 657 910
rect 441 905 442 909
rect 446 905 657 909
rect 441 904 447 905
rect 1108 894 1114 895
rect 1108 890 1109 894
rect 1113 890 1114 894
rect 1108 889 1114 890
rect 693 868 733 869
rect 693 864 727 868
rect 692 863 699 864
rect 692 858 693 863
rect 698 858 699 863
rect 726 863 727 864
rect 732 863 733 868
rect 765 868 801 873
rect 726 862 733 863
rect 750 863 757 864
rect 692 857 699 858
rect 703 859 710 860
rect 703 854 704 859
rect 709 854 710 859
rect 750 858 751 863
rect 756 858 757 863
rect 765 862 766 868
rect 771 867 801 868
rect 771 862 772 867
rect 796 864 801 867
rect 765 861 772 862
rect 795 863 802 864
rect 795 858 796 863
rect 801 858 802 863
rect 824 862 831 863
rect 750 857 757 858
rect 779 857 786 858
rect 795 857 802 858
rect 808 857 814 858
rect 751 854 756 857
rect 703 849 756 854
rect 779 852 780 857
rect 785 852 786 857
rect 808 852 809 857
rect 813 852 814 857
rect 779 851 814 852
rect 780 847 814 851
rect 824 857 825 862
rect 830 857 831 862
rect 906 862 913 863
rect 906 857 907 862
rect 912 857 913 862
rect 991 862 998 863
rect 991 857 992 862
rect 997 857 998 862
rect 824 856 831 857
rect 850 856 857 857
rect 906 856 913 857
rect 931 856 938 857
rect 991 856 998 857
rect 824 851 851 856
rect 856 851 857 856
rect 907 851 932 856
rect 937 851 938 856
rect 824 830 829 851
rect 850 850 857 851
rect 931 850 938 851
rect 988 851 997 856
rect 657 824 829 830
rect 440 806 446 807
rect 440 802 441 806
rect 445 802 578 806
rect 657 804 662 824
rect 440 801 578 802
rect 184 406 190 407
rect 184 402 185 406
rect 189 402 190 406
rect 184 401 190 402
rect 573 42 578 801
rect 656 803 663 804
rect 656 798 657 803
rect 662 798 663 803
rect 656 797 663 798
rect 703 800 756 805
rect 780 803 814 807
rect 692 796 699 797
rect 692 791 693 796
rect 698 791 699 796
rect 703 795 704 800
rect 709 795 710 800
rect 751 797 756 800
rect 779 802 814 803
rect 779 797 780 802
rect 785 797 786 802
rect 808 797 809 802
rect 813 797 814 802
rect 703 794 710 795
rect 750 796 757 797
rect 779 796 786 797
rect 795 796 802 797
rect 808 796 814 797
rect 824 797 831 798
rect 850 797 857 798
rect 930 797 937 798
rect 692 790 699 791
rect 726 791 733 792
rect 726 790 727 791
rect 693 786 727 790
rect 732 786 733 791
rect 750 791 751 796
rect 756 791 757 796
rect 750 790 757 791
rect 765 792 772 793
rect 693 785 733 786
rect 765 786 766 792
rect 771 787 772 792
rect 795 791 796 796
rect 801 791 802 796
rect 824 792 825 797
rect 830 792 851 797
rect 856 792 857 797
rect 824 791 831 792
rect 850 791 857 792
rect 907 792 931 797
rect 936 792 937 797
rect 795 790 802 791
rect 796 787 801 790
rect 771 786 801 787
rect 765 781 801 786
rect 825 764 830 791
rect 656 758 830 764
rect 656 735 661 758
rect 693 736 733 737
rect 655 734 662 735
rect 655 729 656 734
rect 661 729 662 734
rect 693 732 727 736
rect 655 728 662 729
rect 692 731 699 732
rect 692 726 693 731
rect 698 726 699 731
rect 726 731 727 732
rect 732 731 733 736
rect 765 736 801 741
rect 907 739 912 792
rect 930 791 937 792
rect 988 763 993 851
rect 950 758 993 763
rect 726 730 733 731
rect 750 731 757 732
rect 692 725 699 726
rect 703 727 710 728
rect 703 722 704 727
rect 709 722 710 727
rect 750 726 751 731
rect 756 726 757 731
rect 765 730 766 736
rect 771 735 801 736
rect 771 730 772 735
rect 796 732 801 735
rect 906 738 913 739
rect 906 733 907 738
rect 912 733 913 738
rect 906 732 913 733
rect 765 729 772 730
rect 795 731 802 732
rect 795 726 796 731
rect 801 726 802 731
rect 824 730 831 731
rect 750 725 757 726
rect 779 725 786 726
rect 795 725 802 726
rect 808 725 814 726
rect 751 722 756 725
rect 703 717 756 722
rect 779 720 780 725
rect 785 720 786 725
rect 808 720 809 725
rect 813 720 814 725
rect 779 719 814 720
rect 780 715 814 719
rect 824 725 825 730
rect 830 725 831 730
rect 950 725 955 758
rect 1013 735 1020 736
rect 1013 730 1014 735
rect 1019 730 1020 735
rect 1013 729 1020 730
rect 824 724 831 725
rect 850 724 857 725
rect 824 719 851 724
rect 856 719 857 724
rect 950 724 962 725
rect 950 719 956 724
rect 961 719 962 724
rect 824 698 829 719
rect 850 718 857 719
rect 955 718 962 719
rect 657 692 829 698
rect 657 672 662 692
rect 656 671 663 672
rect 656 666 657 671
rect 662 666 663 671
rect 656 665 663 666
rect 703 668 756 673
rect 780 671 814 675
rect 692 664 699 665
rect 692 659 693 664
rect 698 659 699 664
rect 703 663 704 668
rect 709 663 710 668
rect 751 665 756 668
rect 779 670 814 671
rect 779 665 780 670
rect 785 665 786 670
rect 808 665 809 670
rect 813 665 814 670
rect 849 666 856 667
rect 955 666 962 667
rect 703 662 710 663
rect 750 664 757 665
rect 779 664 786 665
rect 795 664 802 665
rect 808 664 814 665
rect 824 665 850 666
rect 692 658 699 659
rect 726 659 733 660
rect 726 658 727 659
rect 693 654 727 658
rect 732 654 733 659
rect 750 659 751 664
rect 756 659 757 664
rect 750 658 757 659
rect 765 660 772 661
rect 693 653 733 654
rect 765 654 766 660
rect 771 655 772 660
rect 795 659 796 664
rect 801 659 802 664
rect 795 658 802 659
rect 824 660 825 665
rect 830 661 850 665
rect 855 661 856 666
rect 830 660 831 661
rect 849 660 856 661
rect 951 661 956 666
rect 961 661 962 666
rect 951 660 962 661
rect 824 659 831 660
rect 796 655 801 658
rect 771 654 801 655
rect 765 649 801 654
rect 824 632 829 659
rect 656 626 829 632
rect 951 632 956 660
rect 951 627 994 632
rect 656 603 661 626
rect 693 604 733 605
rect 655 602 662 603
rect 655 597 656 602
rect 661 597 662 602
rect 693 600 727 604
rect 655 596 662 597
rect 692 599 699 600
rect 692 594 693 599
rect 698 594 699 599
rect 726 599 727 600
rect 732 599 733 604
rect 765 604 801 609
rect 989 608 994 627
rect 726 598 733 599
rect 750 599 757 600
rect 692 593 699 594
rect 703 595 710 596
rect 703 590 704 595
rect 709 590 710 595
rect 750 594 751 599
rect 756 594 757 599
rect 765 598 766 604
rect 771 603 801 604
rect 771 598 772 603
rect 796 600 801 603
rect 988 607 995 608
rect 988 602 989 607
rect 994 602 995 607
rect 988 601 995 602
rect 1014 600 1019 729
rect 1022 600 1029 601
rect 765 597 772 598
rect 795 599 802 600
rect 795 594 796 599
rect 801 594 802 599
rect 824 598 831 599
rect 750 593 757 594
rect 779 593 786 594
rect 795 593 802 594
rect 808 593 814 594
rect 751 590 756 593
rect 703 585 756 590
rect 779 588 780 593
rect 785 588 786 593
rect 808 588 809 593
rect 813 588 814 593
rect 779 587 814 588
rect 780 583 814 587
rect 824 593 825 598
rect 830 593 831 598
rect 906 598 913 599
rect 906 593 907 598
rect 912 593 913 598
rect 1002 595 1023 600
rect 1028 595 1029 600
rect 1002 594 1014 595
rect 1022 594 1029 595
rect 824 592 831 593
rect 850 592 857 593
rect 906 592 913 593
rect 931 592 938 593
rect 824 587 851 592
rect 856 587 857 592
rect 907 587 932 592
rect 937 587 938 592
rect 824 566 829 587
rect 850 586 857 587
rect 931 586 938 587
rect 1002 586 1007 594
rect 657 560 829 566
rect 969 565 1007 586
rect 657 540 662 560
rect 656 539 663 540
rect 656 534 657 539
rect 662 534 663 539
rect 656 533 663 534
rect 703 536 756 541
rect 780 539 814 543
rect 692 532 699 533
rect 692 527 693 532
rect 698 527 699 532
rect 703 531 704 536
rect 709 531 710 536
rect 751 533 756 536
rect 779 538 814 539
rect 779 533 780 538
rect 785 533 786 538
rect 808 533 809 538
rect 813 533 814 538
rect 703 530 710 531
rect 750 532 757 533
rect 779 532 786 533
rect 795 532 802 533
rect 808 532 814 533
rect 824 533 831 534
rect 692 526 699 527
rect 726 527 733 528
rect 726 526 727 527
rect 693 522 727 526
rect 732 522 733 527
rect 750 527 751 532
rect 756 527 757 532
rect 750 526 757 527
rect 765 528 772 529
rect 693 521 733 522
rect 765 522 766 528
rect 771 523 772 528
rect 795 527 796 532
rect 801 527 802 532
rect 824 528 825 533
rect 830 531 831 533
rect 850 531 857 532
rect 930 531 937 532
rect 830 528 851 531
rect 824 527 851 528
rect 795 526 802 527
rect 825 526 851 527
rect 856 526 857 531
rect 796 523 801 526
rect 771 522 801 523
rect 765 517 801 522
rect 825 500 830 526
rect 850 525 857 526
rect 907 526 931 531
rect 936 526 937 531
rect 656 494 830 500
rect 656 471 661 494
rect 693 472 733 473
rect 655 470 662 471
rect 655 465 656 470
rect 661 465 662 470
rect 693 468 727 472
rect 655 464 662 465
rect 692 467 699 468
rect 692 462 693 467
rect 698 462 699 467
rect 726 467 727 468
rect 732 467 733 472
rect 765 472 801 477
rect 907 475 912 526
rect 930 525 937 526
rect 726 466 733 467
rect 750 467 757 468
rect 692 461 699 462
rect 703 463 710 464
rect 703 458 704 463
rect 709 458 710 463
rect 750 462 751 467
rect 756 462 757 467
rect 765 466 766 472
rect 771 471 801 472
rect 771 466 772 471
rect 796 468 801 471
rect 906 474 913 475
rect 906 469 907 474
rect 912 469 913 474
rect 906 468 913 469
rect 765 465 772 466
rect 795 467 802 468
rect 795 462 796 467
rect 801 462 802 467
rect 824 466 831 467
rect 750 461 757 462
rect 779 461 786 462
rect 795 461 802 462
rect 808 461 814 462
rect 751 458 756 461
rect 703 453 756 458
rect 779 456 780 461
rect 785 456 786 461
rect 808 456 809 461
rect 813 456 814 461
rect 779 455 814 456
rect 780 451 814 455
rect 824 461 825 466
rect 830 461 831 466
rect 824 460 831 461
rect 850 460 857 461
rect 824 455 851 460
rect 856 455 857 460
rect 969 456 974 565
rect 1019 527 1026 528
rect 1019 522 1020 527
rect 1025 522 1026 527
rect 1019 521 1026 522
rect 926 455 974 456
rect 824 434 829 455
rect 850 454 857 455
rect 657 428 829 434
rect 895 450 974 455
rect 1020 459 1025 521
rect 1020 453 1087 459
rect 657 408 662 428
rect 656 407 663 408
rect 656 402 657 407
rect 662 402 663 407
rect 656 401 663 402
rect 703 404 756 409
rect 780 407 814 411
rect 895 407 900 450
rect 692 400 699 401
rect 692 395 693 400
rect 698 395 699 400
rect 703 399 704 404
rect 709 399 710 404
rect 751 401 756 404
rect 779 406 814 407
rect 779 401 780 406
rect 785 401 786 406
rect 808 401 809 406
rect 813 401 814 406
rect 894 406 901 407
rect 703 398 710 399
rect 750 400 757 401
rect 779 400 786 401
rect 795 400 802 401
rect 808 400 814 401
rect 824 401 831 402
rect 692 394 699 395
rect 726 395 733 396
rect 726 394 727 395
rect 693 390 727 394
rect 732 390 733 395
rect 750 395 751 400
rect 756 395 757 400
rect 750 394 757 395
rect 765 396 772 397
rect 693 389 733 390
rect 765 390 766 396
rect 771 391 772 396
rect 795 395 796 400
rect 801 395 802 400
rect 824 396 825 401
rect 830 396 831 401
rect 894 401 895 406
rect 900 401 901 406
rect 964 404 1017 409
rect 1041 407 1075 411
rect 1082 407 1087 453
rect 894 400 901 401
rect 953 400 960 401
rect 824 395 831 396
rect 849 395 856 396
rect 795 394 802 395
rect 796 391 801 394
rect 771 390 801 391
rect 826 390 850 395
rect 855 390 856 395
rect 953 395 954 400
rect 959 395 960 400
rect 964 399 965 404
rect 970 399 971 404
rect 1012 401 1017 404
rect 1040 406 1075 407
rect 1040 401 1041 406
rect 1046 401 1047 406
rect 1069 401 1070 406
rect 1074 401 1075 406
rect 964 398 971 399
rect 1011 400 1018 401
rect 1040 400 1047 401
rect 1056 400 1063 401
rect 1069 400 1075 401
rect 1081 406 1088 407
rect 1081 401 1082 406
rect 1087 401 1088 406
rect 1081 400 1088 401
rect 953 394 960 395
rect 987 395 994 396
rect 987 394 988 395
rect 765 385 801 390
rect 849 389 856 390
rect 954 390 988 394
rect 993 390 994 395
rect 1011 395 1012 400
rect 1017 395 1018 400
rect 1011 394 1018 395
rect 1026 396 1033 397
rect 954 389 994 390
rect 1026 390 1027 396
rect 1032 391 1033 396
rect 1056 395 1057 400
rect 1062 395 1063 400
rect 1056 394 1063 395
rect 1057 391 1062 394
rect 1032 390 1062 391
rect 1026 385 1062 390
rect 1109 362 1114 889
rect 956 357 1114 362
rect 956 297 961 357
rect 955 296 961 297
rect 955 292 956 296
rect 960 292 961 296
rect 955 291 961 292
rect 1081 229 1115 234
rect 1081 215 1086 229
rect 1080 214 1086 215
rect 1080 210 1081 214
rect 1085 210 1086 214
rect 1080 209 1086 210
rect 573 41 579 42
rect 573 37 574 41
rect 578 37 579 41
rect 573 36 579 37
rect 185 0 1115 5
<< labels >>
rlabel metal2 596 984 596 984 1 GND!
rlabel metal2 584 984 584 984 1 Vdd!
rlabel metal2 609 983 609 983 4 f_clk_b
rlabel metal2 621 982 621 982 5 f_clk
rlabel metal2 645 983 645 983 5 p_clk
rlabel metal2 633 983 633 983 5 p_clk_b
rlabel metal2 433 972 437 994 1 fin2
rlabel metal2 316 973 320 995 1 fin1
rlabel metal2 618 955 624 964 1 f_clk
rlabel metal2 606 956 612 965 1 f_clk_b
rlabel metal2 786 899 794 900 1 s0
rlabel metal2 915 899 917 901 1 s1
rlabel metal2 983 898 985 900 1 s2
rlabel metal2 1179 896 1181 898 7 s3
rlabel m3contact 1015 730 1017 732 1 out
rlabel metal1 656 857 659 859 1 fin
<< end >>
