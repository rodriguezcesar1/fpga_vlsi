magic
tech scmos
timestamp 1607526808
<< ntransistor >>
rect 425 294 427 298
rect 441 294 443 298
rect 460 294 462 298
rect 480 294 482 298
rect 485 294 487 298
rect 511 294 513 298
rect 536 294 538 298
rect 556 294 558 298
rect 561 294 563 298
rect 590 294 592 298
rect 611 294 613 298
<< ptransistor >>
rect 425 313 427 321
rect 441 313 443 321
rect 460 314 462 322
rect 480 313 482 321
rect 485 313 487 321
rect 511 313 513 321
rect 536 314 538 322
rect 556 313 558 321
rect 561 313 563 321
rect 590 313 592 321
rect 611 313 613 321
<< ndiffusion >>
rect 424 294 425 298
rect 427 294 428 298
rect 440 294 441 298
rect 443 294 444 298
rect 459 294 460 298
rect 462 294 463 298
rect 475 294 480 298
rect 482 294 485 298
rect 487 294 488 298
rect 510 294 511 298
rect 513 294 514 298
rect 535 294 536 298
rect 538 294 539 298
rect 551 294 556 298
rect 558 294 561 298
rect 563 294 564 298
rect 589 294 590 298
rect 592 294 593 298
rect 610 294 611 298
rect 613 294 614 298
<< pdiffusion >>
rect 424 313 425 321
rect 427 313 428 321
rect 440 313 441 321
rect 443 313 444 321
rect 459 314 460 322
rect 462 314 463 322
rect 475 313 480 321
rect 482 313 485 321
rect 487 313 488 321
rect 510 313 511 321
rect 513 313 514 321
rect 535 314 536 322
rect 538 314 539 322
rect 551 313 556 321
rect 558 313 561 321
rect 563 313 564 321
rect 589 313 590 321
rect 592 313 593 321
rect 610 313 611 321
rect 613 313 614 321
<< ndcontact >>
rect 420 294 424 298
rect 428 294 432 298
rect 436 294 440 298
rect 444 294 448 298
rect 455 294 459 298
rect 463 294 467 298
rect 471 294 475 298
rect 488 294 492 298
rect 506 294 510 298
rect 514 294 518 298
rect 531 294 535 298
rect 539 294 543 298
rect 547 294 551 298
rect 564 294 568 298
rect 585 294 589 298
rect 593 294 597 298
rect 606 294 610 298
rect 614 294 618 298
<< pdcontact >>
rect 420 313 424 321
rect 428 313 432 321
rect 436 313 440 321
rect 444 313 448 321
rect 455 314 459 322
rect 463 314 467 322
rect 471 313 475 321
rect 488 313 492 321
rect 506 313 510 321
rect 514 313 518 321
rect 531 314 535 322
rect 539 314 543 322
rect 547 313 551 321
rect 564 313 568 321
rect 585 313 589 321
rect 593 313 597 321
rect 606 313 610 321
rect 614 313 618 321
<< psubstratepcontact >>
rect 413 278 417 282
rect 431 278 435 282
rect 451 278 455 282
rect 464 278 468 282
rect 501 278 505 282
rect 523 278 527 282
rect 540 278 544 282
rect 575 278 579 282
<< nsubstratencontact >>
rect 413 331 417 335
rect 431 331 435 335
rect 451 331 455 335
rect 464 331 468 335
rect 501 331 505 335
rect 523 331 527 335
rect 540 331 544 335
rect 575 331 579 335
<< polysilicon >>
rect 441 328 443 331
rect 485 328 487 331
rect 511 328 513 331
rect 561 328 563 331
rect 441 324 442 328
rect 511 324 512 328
rect 425 321 427 323
rect 441 321 443 324
rect 460 322 462 324
rect 480 321 482 323
rect 485 321 487 324
rect 511 321 513 324
rect 536 322 538 324
rect 425 298 427 313
rect 441 311 443 313
rect 441 298 443 300
rect 460 298 462 314
rect 556 321 558 323
rect 561 321 563 324
rect 590 321 592 323
rect 611 321 613 323
rect 480 307 482 313
rect 485 311 487 313
rect 511 311 513 313
rect 476 303 482 307
rect 480 298 482 303
rect 485 298 487 300
rect 511 298 513 300
rect 536 298 538 314
rect 556 307 558 313
rect 561 311 563 313
rect 552 303 558 307
rect 556 298 558 303
rect 561 298 563 300
rect 590 298 592 313
rect 611 298 613 313
rect 425 292 427 294
rect 441 290 443 294
rect 460 292 462 294
rect 480 292 482 294
rect 442 286 443 290
rect 485 289 487 294
rect 511 290 513 294
rect 536 292 538 294
rect 556 292 558 294
rect 441 283 443 286
rect 486 285 487 289
rect 512 286 513 290
rect 561 289 563 294
rect 590 292 592 294
rect 611 292 613 294
rect 485 283 487 285
rect 511 282 513 286
rect 562 285 563 289
rect 561 283 563 285
<< polycontact >>
rect 442 324 446 328
rect 485 324 489 328
rect 512 324 516 328
rect 561 324 565 328
rect 421 303 425 307
rect 456 304 460 308
rect 472 303 476 307
rect 532 304 536 308
rect 548 303 552 307
rect 586 303 590 307
rect 607 303 611 307
rect 438 286 442 290
rect 482 285 486 289
rect 508 286 512 290
rect 558 285 562 289
<< metal1 >>
rect 413 340 447 344
rect 451 340 474 344
rect 478 340 503 344
rect 507 340 550 344
rect 554 340 618 344
rect 417 331 431 335
rect 435 331 451 335
rect 455 331 464 335
rect 468 331 501 335
rect 505 331 523 335
rect 527 331 540 335
rect 544 331 575 335
rect 579 331 618 335
rect 420 321 423 331
rect 446 324 447 328
rect 455 322 458 331
rect 416 303 421 306
rect 429 306 432 313
rect 436 306 439 313
rect 429 303 439 306
rect 429 298 432 303
rect 436 298 439 303
rect 445 308 448 313
rect 445 307 450 308
rect 445 304 456 307
rect 464 306 467 314
rect 471 321 474 331
rect 489 324 496 328
rect 516 324 517 328
rect 531 322 534 331
rect 489 307 492 313
rect 445 298 448 304
rect 464 303 472 306
rect 488 306 492 307
rect 506 306 509 313
rect 488 303 509 306
rect 464 298 467 303
rect 489 298 492 303
rect 506 298 509 303
rect 515 307 518 313
rect 524 307 528 308
rect 515 304 532 307
rect 540 306 543 314
rect 547 321 550 331
rect 565 324 571 328
rect 585 321 588 331
rect 606 321 609 331
rect 565 307 568 313
rect 515 298 518 304
rect 540 303 548 306
rect 564 306 568 307
rect 580 306 583 307
rect 564 303 586 306
rect 540 298 543 303
rect 565 298 568 303
rect 579 302 585 303
rect 594 298 597 313
rect 601 306 604 307
rect 600 303 607 306
rect 600 302 606 303
rect 615 298 618 313
rect 420 282 423 294
rect 437 286 438 290
rect 455 282 458 294
rect 471 282 474 294
rect 481 285 482 289
rect 507 286 508 290
rect 531 282 534 294
rect 547 282 550 294
rect 557 285 558 289
rect 585 282 588 294
rect 606 282 609 294
rect 417 278 431 282
rect 435 278 451 282
rect 455 278 464 282
rect 468 278 501 282
rect 505 278 523 282
rect 527 278 540 282
rect 544 278 575 282
rect 579 278 618 282
rect 413 270 433 274
rect 437 270 497 274
rect 501 270 518 274
rect 522 270 572 274
rect 576 270 618 274
<< m2contact >>
rect 447 340 451 344
rect 474 340 478 344
rect 503 340 507 344
rect 550 340 554 344
rect 447 324 451 328
rect 496 324 500 328
rect 517 324 521 328
rect 571 324 575 328
rect 433 286 437 290
rect 477 285 481 289
rect 503 286 507 290
rect 553 285 557 289
rect 433 270 437 274
rect 497 270 501 274
rect 518 270 522 274
rect 572 270 576 274
<< metal2 >>
rect 447 328 451 340
rect 451 304 452 307
rect 433 274 437 286
rect 474 285 477 340
rect 497 274 500 324
rect 503 290 506 340
rect 518 274 521 324
rect 550 285 553 340
rect 572 274 575 324
rect 578 303 579 306
<< m3contact >>
rect 446 304 451 309
rect 488 303 493 308
rect 524 304 529 309
rect 564 303 569 308
rect 579 302 584 307
rect 600 302 605 307
<< metal3 >>
rect 524 313 605 318
rect 524 310 529 313
rect 445 309 452 310
rect 523 309 530 310
rect 445 304 446 309
rect 451 308 494 309
rect 451 304 488 308
rect 445 303 452 304
rect 487 303 488 304
rect 493 303 494 308
rect 523 304 524 309
rect 529 308 570 309
rect 600 308 605 313
rect 529 304 564 308
rect 523 303 530 304
rect 563 303 564 304
rect 569 303 570 308
rect 487 302 494 303
rect 524 297 529 303
rect 563 302 570 303
rect 578 307 585 308
rect 578 302 579 307
rect 584 302 585 307
rect 578 301 585 302
rect 599 307 606 308
rect 599 302 600 307
rect 605 302 606 307
rect 599 301 606 302
rect 579 297 584 301
rect 524 292 584 297
<< labels >>
rlabel metal1 416 303 420 306 1 D
rlabel metal1 615 301 618 308 7 Q
rlabel metal1 594 301 597 308 1 ~Q
<< end >>
