magic
tech scmos
timestamp 1607527890
<< ntransistor >>
rect 12 24 14 28
rect 28 24 30 28
rect 47 24 49 28
rect 67 24 69 28
rect 72 24 74 28
rect 98 24 100 28
rect 123 24 125 28
rect 143 24 145 28
rect 148 24 150 28
rect 177 24 179 28
rect 198 24 200 28
rect 214 24 216 28
rect 230 24 232 28
rect 249 24 251 28
rect 269 24 271 28
rect 274 24 276 28
rect 300 24 302 28
rect 325 24 327 28
rect 345 24 347 28
rect 350 24 352 28
rect 379 24 381 28
rect 400 24 402 28
rect 416 24 418 28
rect 432 24 434 28
rect 451 24 453 28
rect 471 24 473 28
rect 476 24 478 28
rect 502 24 504 28
rect 527 24 529 28
rect 547 24 549 28
rect 552 24 554 28
rect 581 24 583 28
rect 602 24 604 28
rect 618 24 620 28
rect 634 24 636 28
rect 653 24 655 28
rect 673 24 675 28
rect 678 24 680 28
rect 704 24 706 28
rect 729 24 731 28
rect 749 24 751 28
rect 754 24 756 28
rect 783 24 785 28
rect 804 24 806 28
<< ptransistor >>
rect 12 43 14 51
rect 28 43 30 51
rect 47 44 49 52
rect 67 43 69 51
rect 72 43 74 51
rect 98 43 100 51
rect 123 44 125 52
rect 143 43 145 51
rect 148 43 150 51
rect 177 43 179 51
rect 198 43 200 51
rect 214 43 216 51
rect 230 43 232 51
rect 249 44 251 52
rect 269 43 271 51
rect 274 43 276 51
rect 300 43 302 51
rect 325 44 327 52
rect 345 43 347 51
rect 350 43 352 51
rect 379 43 381 51
rect 400 43 402 51
rect 416 43 418 51
rect 432 43 434 51
rect 451 44 453 52
rect 471 43 473 51
rect 476 43 478 51
rect 502 43 504 51
rect 527 44 529 52
rect 547 43 549 51
rect 552 43 554 51
rect 581 43 583 51
rect 602 43 604 51
rect 618 43 620 51
rect 634 43 636 51
rect 653 44 655 52
rect 673 43 675 51
rect 678 43 680 51
rect 704 43 706 51
rect 729 44 731 52
rect 749 43 751 51
rect 754 43 756 51
rect 783 43 785 51
rect 804 43 806 51
<< ndiffusion >>
rect 11 24 12 28
rect 14 24 15 28
rect 27 24 28 28
rect 30 24 31 28
rect 46 24 47 28
rect 49 24 50 28
rect 62 24 67 28
rect 69 24 72 28
rect 74 24 75 28
rect 97 24 98 28
rect 100 24 101 28
rect 122 24 123 28
rect 125 24 126 28
rect 138 24 143 28
rect 145 24 148 28
rect 150 24 151 28
rect 176 24 177 28
rect 179 24 180 28
rect 197 24 198 28
rect 200 24 201 28
rect 213 24 214 28
rect 216 24 217 28
rect 229 24 230 28
rect 232 24 233 28
rect 248 24 249 28
rect 251 24 252 28
rect 264 24 269 28
rect 271 24 274 28
rect 276 24 277 28
rect 299 24 300 28
rect 302 24 303 28
rect 324 24 325 28
rect 327 24 328 28
rect 340 24 345 28
rect 347 24 350 28
rect 352 24 353 28
rect 378 24 379 28
rect 381 24 382 28
rect 399 24 400 28
rect 402 24 403 28
rect 415 24 416 28
rect 418 24 419 28
rect 431 24 432 28
rect 434 24 435 28
rect 450 24 451 28
rect 453 24 454 28
rect 466 24 471 28
rect 473 24 476 28
rect 478 24 479 28
rect 501 24 502 28
rect 504 24 505 28
rect 526 24 527 28
rect 529 24 530 28
rect 542 24 547 28
rect 549 24 552 28
rect 554 24 555 28
rect 580 24 581 28
rect 583 24 584 28
rect 601 24 602 28
rect 604 24 605 28
rect 617 24 618 28
rect 620 24 621 28
rect 633 24 634 28
rect 636 24 637 28
rect 652 24 653 28
rect 655 24 656 28
rect 668 24 673 28
rect 675 24 678 28
rect 680 24 681 28
rect 703 24 704 28
rect 706 24 707 28
rect 728 24 729 28
rect 731 24 732 28
rect 744 24 749 28
rect 751 24 754 28
rect 756 24 757 28
rect 782 24 783 28
rect 785 24 786 28
rect 803 24 804 28
rect 806 24 807 28
<< pdiffusion >>
rect 11 43 12 51
rect 14 43 15 51
rect 27 43 28 51
rect 30 43 31 51
rect 46 44 47 52
rect 49 44 50 52
rect 62 43 67 51
rect 69 43 72 51
rect 74 43 75 51
rect 97 43 98 51
rect 100 43 101 51
rect 122 44 123 52
rect 125 44 126 52
rect 138 43 143 51
rect 145 43 148 51
rect 150 43 151 51
rect 176 43 177 51
rect 179 43 180 51
rect 197 43 198 51
rect 200 43 201 51
rect 213 43 214 51
rect 216 43 217 51
rect 229 43 230 51
rect 232 43 233 51
rect 248 44 249 52
rect 251 44 252 52
rect 264 43 269 51
rect 271 43 274 51
rect 276 43 277 51
rect 299 43 300 51
rect 302 43 303 51
rect 324 44 325 52
rect 327 44 328 52
rect 340 43 345 51
rect 347 43 350 51
rect 352 43 353 51
rect 378 43 379 51
rect 381 43 382 51
rect 399 43 400 51
rect 402 43 403 51
rect 415 43 416 51
rect 418 43 419 51
rect 431 43 432 51
rect 434 43 435 51
rect 450 44 451 52
rect 453 44 454 52
rect 466 43 471 51
rect 473 43 476 51
rect 478 43 479 51
rect 501 43 502 51
rect 504 43 505 51
rect 526 44 527 52
rect 529 44 530 52
rect 542 43 547 51
rect 549 43 552 51
rect 554 43 555 51
rect 580 43 581 51
rect 583 43 584 51
rect 601 43 602 51
rect 604 43 605 51
rect 617 43 618 51
rect 620 43 621 51
rect 633 43 634 51
rect 636 43 637 51
rect 652 44 653 52
rect 655 44 656 52
rect 668 43 673 51
rect 675 43 678 51
rect 680 43 681 51
rect 703 43 704 51
rect 706 43 707 51
rect 728 44 729 52
rect 731 44 732 52
rect 744 43 749 51
rect 751 43 754 51
rect 756 43 757 51
rect 782 43 783 51
rect 785 43 786 51
rect 803 43 804 51
rect 806 43 807 51
<< ndcontact >>
rect 7 24 11 28
rect 15 24 19 28
rect 23 24 27 28
rect 31 24 35 28
rect 42 24 46 28
rect 50 24 54 28
rect 58 24 62 28
rect 75 24 79 28
rect 93 24 97 28
rect 101 24 105 28
rect 118 24 122 28
rect 126 24 130 28
rect 134 24 138 28
rect 151 24 155 28
rect 172 24 176 28
rect 180 24 184 28
rect 193 24 197 28
rect 201 24 205 28
rect 209 24 213 28
rect 217 24 221 28
rect 225 24 229 28
rect 233 24 237 28
rect 244 24 248 28
rect 252 24 256 28
rect 260 24 264 28
rect 277 24 281 28
rect 295 24 299 28
rect 303 24 307 28
rect 320 24 324 28
rect 328 24 332 28
rect 336 24 340 28
rect 353 24 357 28
rect 374 24 378 28
rect 382 24 386 28
rect 395 24 399 28
rect 403 24 407 28
rect 411 24 415 28
rect 419 24 423 28
rect 427 24 431 28
rect 435 24 439 28
rect 446 24 450 28
rect 454 24 458 28
rect 462 24 466 28
rect 479 24 483 28
rect 497 24 501 28
rect 505 24 509 28
rect 522 24 526 28
rect 530 24 534 28
rect 538 24 542 28
rect 555 24 559 28
rect 576 24 580 28
rect 584 24 588 28
rect 597 24 601 28
rect 605 24 609 28
rect 613 24 617 28
rect 621 24 625 28
rect 629 24 633 28
rect 637 24 641 28
rect 648 24 652 28
rect 656 24 660 28
rect 664 24 668 28
rect 681 24 685 28
rect 699 24 703 28
rect 707 24 711 28
rect 724 24 728 28
rect 732 24 736 28
rect 740 24 744 28
rect 757 24 761 28
rect 778 24 782 28
rect 786 24 790 28
rect 799 24 803 28
rect 807 24 811 28
<< pdcontact >>
rect 7 43 11 51
rect 15 43 19 51
rect 23 43 27 51
rect 31 43 35 51
rect 42 44 46 52
rect 50 44 54 52
rect 58 43 62 51
rect 75 43 79 51
rect 93 43 97 51
rect 101 43 105 51
rect 118 44 122 52
rect 126 44 130 52
rect 134 43 138 51
rect 151 43 155 51
rect 172 43 176 51
rect 180 43 184 51
rect 193 43 197 51
rect 201 43 205 51
rect 209 43 213 51
rect 217 43 221 51
rect 225 43 229 51
rect 233 43 237 51
rect 244 44 248 52
rect 252 44 256 52
rect 260 43 264 51
rect 277 43 281 51
rect 295 43 299 51
rect 303 43 307 51
rect 320 44 324 52
rect 328 44 332 52
rect 336 43 340 51
rect 353 43 357 51
rect 374 43 378 51
rect 382 43 386 51
rect 395 43 399 51
rect 403 43 407 51
rect 411 43 415 51
rect 419 43 423 51
rect 427 43 431 51
rect 435 43 439 51
rect 446 44 450 52
rect 454 44 458 52
rect 462 43 466 51
rect 479 43 483 51
rect 497 43 501 51
rect 505 43 509 51
rect 522 44 526 52
rect 530 44 534 52
rect 538 43 542 51
rect 555 43 559 51
rect 576 43 580 51
rect 584 43 588 51
rect 597 43 601 51
rect 605 43 609 51
rect 613 43 617 51
rect 621 43 625 51
rect 629 43 633 51
rect 637 43 641 51
rect 648 44 652 52
rect 656 44 660 52
rect 664 43 668 51
rect 681 43 685 51
rect 699 43 703 51
rect 707 43 711 51
rect 724 44 728 52
rect 732 44 736 52
rect 740 43 744 51
rect 757 43 761 51
rect 778 43 782 51
rect 786 43 790 51
rect 799 43 803 51
rect 807 43 811 51
<< psubstratepcontact >>
rect 0 8 4 12
rect 18 8 22 12
rect 38 8 42 12
rect 51 8 55 12
rect 88 8 92 12
rect 110 8 114 12
rect 127 8 131 12
rect 162 8 166 12
rect 205 8 209 12
rect 220 8 224 12
rect 240 8 244 12
rect 253 8 257 12
rect 290 8 294 12
rect 312 8 316 12
rect 329 8 333 12
rect 364 8 368 12
rect 407 8 411 12
rect 422 8 426 12
rect 442 8 446 12
rect 455 8 459 12
rect 492 8 496 12
rect 514 8 518 12
rect 531 8 535 12
rect 566 8 570 12
rect 609 8 613 12
rect 624 8 628 12
rect 644 8 648 12
rect 657 8 661 12
rect 694 8 698 12
rect 716 8 720 12
rect 733 8 737 12
rect 768 8 772 12
<< nsubstratencontact >>
rect 0 61 4 65
rect 18 61 22 65
rect 38 61 42 65
rect 51 61 55 65
rect 88 61 92 65
rect 110 61 114 65
rect 127 61 131 65
rect 162 61 166 65
rect 205 61 209 65
rect 220 61 224 65
rect 240 61 244 65
rect 253 61 257 65
rect 290 61 294 65
rect 312 61 316 65
rect 329 61 333 65
rect 364 61 368 65
rect 407 61 411 65
rect 422 61 426 65
rect 442 61 446 65
rect 455 61 459 65
rect 492 61 496 65
rect 514 61 518 65
rect 531 61 535 65
rect 566 61 570 65
rect 609 61 613 65
rect 624 61 628 65
rect 644 61 648 65
rect 657 61 661 65
rect 694 61 698 65
rect 716 61 720 65
rect 733 61 737 65
rect 768 61 772 65
<< polysilicon >>
rect 28 58 30 61
rect 72 58 74 61
rect 98 58 100 61
rect 148 58 150 61
rect 230 58 232 61
rect 274 58 276 61
rect 300 58 302 61
rect 350 58 352 61
rect 432 58 434 61
rect 476 58 478 61
rect 502 58 504 61
rect 552 58 554 61
rect 634 58 636 61
rect 678 58 680 61
rect 704 58 706 61
rect 754 58 756 61
rect 28 54 29 58
rect 98 54 99 58
rect 230 54 231 58
rect 300 54 301 58
rect 432 54 433 58
rect 502 54 503 58
rect 634 54 635 58
rect 704 54 705 58
rect 12 51 14 53
rect 28 51 30 54
rect 47 52 49 54
rect 67 51 69 53
rect 72 51 74 54
rect 98 51 100 54
rect 123 52 125 54
rect 12 28 14 43
rect 28 41 30 43
rect 28 28 30 30
rect 47 28 49 44
rect 143 51 145 53
rect 148 51 150 54
rect 177 51 179 53
rect 198 51 200 53
rect 214 51 216 53
rect 230 51 232 54
rect 249 52 251 54
rect 67 37 69 43
rect 72 41 74 43
rect 98 41 100 43
rect 63 33 69 37
rect 67 28 69 33
rect 72 28 74 30
rect 98 28 100 30
rect 123 28 125 44
rect 269 51 271 53
rect 274 51 276 54
rect 300 51 302 54
rect 325 52 327 54
rect 143 37 145 43
rect 148 41 150 43
rect 139 33 145 37
rect 143 28 145 33
rect 148 28 150 30
rect 177 28 179 43
rect 198 28 200 43
rect 214 28 216 43
rect 230 41 232 43
rect 230 28 232 30
rect 249 28 251 44
rect 345 51 347 53
rect 350 51 352 54
rect 379 51 381 53
rect 400 51 402 53
rect 416 51 418 53
rect 432 51 434 54
rect 451 52 453 54
rect 269 37 271 43
rect 274 41 276 43
rect 300 41 302 43
rect 265 33 271 37
rect 269 28 271 33
rect 274 28 276 30
rect 300 28 302 30
rect 325 28 327 44
rect 471 51 473 53
rect 476 51 478 54
rect 502 51 504 54
rect 527 52 529 54
rect 345 37 347 43
rect 350 41 352 43
rect 341 33 347 37
rect 345 28 347 33
rect 350 28 352 30
rect 379 28 381 43
rect 400 28 402 43
rect 416 28 418 43
rect 432 41 434 43
rect 432 28 434 30
rect 451 28 453 44
rect 547 51 549 53
rect 552 51 554 54
rect 581 51 583 53
rect 602 51 604 53
rect 618 51 620 53
rect 634 51 636 54
rect 653 52 655 54
rect 471 37 473 43
rect 476 41 478 43
rect 502 41 504 43
rect 467 33 473 37
rect 471 28 473 33
rect 476 28 478 30
rect 502 28 504 30
rect 527 28 529 44
rect 673 51 675 53
rect 678 51 680 54
rect 704 51 706 54
rect 729 52 731 54
rect 547 37 549 43
rect 552 41 554 43
rect 543 33 549 37
rect 547 28 549 33
rect 552 28 554 30
rect 581 28 583 43
rect 602 28 604 43
rect 618 28 620 43
rect 634 41 636 43
rect 634 28 636 30
rect 653 28 655 44
rect 749 51 751 53
rect 754 51 756 54
rect 783 51 785 53
rect 804 51 806 53
rect 673 37 675 43
rect 678 41 680 43
rect 704 41 706 43
rect 669 33 675 37
rect 673 28 675 33
rect 678 28 680 30
rect 704 28 706 30
rect 729 28 731 44
rect 749 37 751 43
rect 754 41 756 43
rect 745 33 751 37
rect 749 28 751 33
rect 754 28 756 30
rect 783 28 785 43
rect 804 28 806 43
rect 12 22 14 24
rect 28 20 30 24
rect 47 22 49 24
rect 67 22 69 24
rect 29 16 30 20
rect 72 19 74 24
rect 98 20 100 24
rect 123 22 125 24
rect 143 22 145 24
rect 28 13 30 16
rect 73 15 74 19
rect 99 16 100 20
rect 148 19 150 24
rect 177 22 179 24
rect 198 22 200 24
rect 214 22 216 24
rect 230 20 232 24
rect 249 22 251 24
rect 269 22 271 24
rect 72 13 74 15
rect 98 12 100 16
rect 149 15 150 19
rect 231 16 232 20
rect 274 19 276 24
rect 300 20 302 24
rect 325 22 327 24
rect 345 22 347 24
rect 148 13 150 15
rect 230 13 232 16
rect 275 15 276 19
rect 301 16 302 20
rect 350 19 352 24
rect 379 22 381 24
rect 400 22 402 24
rect 416 22 418 24
rect 432 20 434 24
rect 451 22 453 24
rect 471 22 473 24
rect 274 13 276 15
rect 300 12 302 16
rect 351 15 352 19
rect 433 16 434 20
rect 476 19 478 24
rect 502 20 504 24
rect 527 22 529 24
rect 547 22 549 24
rect 350 13 352 15
rect 432 13 434 16
rect 477 15 478 19
rect 503 16 504 20
rect 552 19 554 24
rect 581 22 583 24
rect 602 22 604 24
rect 618 22 620 24
rect 634 20 636 24
rect 653 22 655 24
rect 673 22 675 24
rect 476 13 478 15
rect 502 12 504 16
rect 553 15 554 19
rect 635 16 636 20
rect 678 19 680 24
rect 704 20 706 24
rect 729 22 731 24
rect 749 22 751 24
rect 552 13 554 15
rect 634 13 636 16
rect 679 15 680 19
rect 705 16 706 20
rect 754 19 756 24
rect 783 22 785 24
rect 804 22 806 24
rect 678 13 680 15
rect 704 12 706 16
rect 755 15 756 19
rect 754 13 756 15
<< polycontact >>
rect 29 54 33 58
rect 72 54 76 58
rect 99 54 103 58
rect 148 54 152 58
rect 231 54 235 58
rect 274 54 278 58
rect 301 54 305 58
rect 350 54 354 58
rect 433 54 437 58
rect 476 54 480 58
rect 503 54 507 58
rect 552 54 556 58
rect 635 54 639 58
rect 678 54 682 58
rect 705 54 709 58
rect 754 54 758 58
rect 8 33 12 37
rect 43 34 47 38
rect 59 33 63 37
rect 119 34 123 38
rect 135 33 139 37
rect 173 33 177 37
rect 194 33 198 37
rect 210 33 214 37
rect 245 34 249 38
rect 261 33 265 37
rect 321 34 325 38
rect 337 33 341 37
rect 375 33 379 37
rect 396 33 400 37
rect 412 33 416 37
rect 447 34 451 38
rect 463 33 467 37
rect 523 34 527 38
rect 539 33 543 37
rect 577 33 581 37
rect 598 33 602 37
rect 614 33 618 37
rect 649 34 653 38
rect 665 33 669 37
rect 725 34 729 38
rect 741 33 745 37
rect 779 33 783 37
rect 800 33 804 37
rect 25 16 29 20
rect 69 15 73 19
rect 95 16 99 20
rect 145 15 149 19
rect 227 16 231 20
rect 271 15 275 19
rect 297 16 301 20
rect 347 15 351 19
rect 429 16 433 20
rect 473 15 477 19
rect 499 16 503 20
rect 549 15 553 19
rect 631 16 635 20
rect 675 15 679 19
rect 701 16 705 20
rect 751 15 755 19
<< metal1 >>
rect 0 70 34 74
rect 38 70 61 74
rect 65 70 90 74
rect 94 70 137 74
rect 141 70 236 74
rect 240 70 263 74
rect 267 70 292 74
rect 296 70 339 74
rect 343 70 438 74
rect 442 70 465 74
rect 469 70 494 74
rect 498 70 541 74
rect 545 70 640 74
rect 644 70 667 74
rect 671 70 696 74
rect 700 70 743 74
rect 747 70 811 74
rect 4 61 18 65
rect 22 61 38 65
rect 42 61 51 65
rect 55 61 88 65
rect 92 61 110 65
rect 114 61 127 65
rect 131 61 162 65
rect 166 61 205 65
rect 209 61 220 65
rect 224 61 240 65
rect 244 61 253 65
rect 257 61 290 65
rect 294 61 312 65
rect 316 61 329 65
rect 333 61 364 65
rect 368 61 407 65
rect 411 61 422 65
rect 426 61 442 65
rect 446 61 455 65
rect 459 61 492 65
rect 496 61 514 65
rect 518 61 531 65
rect 535 61 566 65
rect 570 61 609 65
rect 613 61 624 65
rect 628 61 644 65
rect 648 61 657 65
rect 661 61 694 65
rect 698 61 716 65
rect 720 61 733 65
rect 737 61 768 65
rect 772 61 811 65
rect 7 51 10 61
rect 33 54 34 58
rect 42 52 45 61
rect 3 33 8 36
rect 16 36 19 43
rect 23 36 26 43
rect 16 33 26 36
rect 16 28 19 33
rect 23 28 26 33
rect 32 38 35 43
rect 32 37 37 38
rect 32 34 43 37
rect 51 36 54 44
rect 58 51 61 61
rect 76 54 83 58
rect 103 54 104 58
rect 118 52 121 61
rect 76 37 79 43
rect 32 28 35 34
rect 51 33 59 36
rect 75 36 79 37
rect 93 36 96 43
rect 75 33 96 36
rect 51 28 54 33
rect 76 28 79 33
rect 93 28 96 33
rect 102 37 105 43
rect 111 37 115 38
rect 102 34 119 37
rect 127 36 130 44
rect 134 51 137 61
rect 152 54 158 58
rect 172 51 175 61
rect 193 51 196 61
rect 209 51 212 61
rect 235 54 236 58
rect 244 52 247 61
rect 152 37 155 43
rect 102 28 105 34
rect 127 33 135 36
rect 151 36 155 37
rect 167 36 170 37
rect 151 33 173 36
rect 127 28 130 33
rect 152 28 155 33
rect 166 32 172 33
rect 181 28 184 43
rect 188 36 191 37
rect 187 33 194 36
rect 202 36 205 43
rect 202 33 210 36
rect 218 36 221 43
rect 225 36 228 43
rect 218 33 228 36
rect 187 32 193 33
rect 202 28 205 33
rect 218 28 221 33
rect 225 28 228 33
rect 234 38 237 43
rect 234 37 239 38
rect 234 34 245 37
rect 253 36 256 44
rect 260 51 263 61
rect 278 54 285 58
rect 305 54 306 58
rect 320 52 323 61
rect 278 37 281 43
rect 234 28 237 34
rect 253 33 261 36
rect 277 36 281 37
rect 295 36 298 43
rect 277 33 298 36
rect 253 28 256 33
rect 278 28 281 33
rect 295 28 298 33
rect 304 37 307 43
rect 313 37 317 38
rect 304 34 321 37
rect 329 36 332 44
rect 336 51 339 61
rect 354 54 360 58
rect 374 51 377 61
rect 395 51 398 61
rect 411 51 414 61
rect 437 54 438 58
rect 446 52 449 61
rect 354 37 357 43
rect 304 28 307 34
rect 329 33 337 36
rect 353 36 357 37
rect 369 36 372 37
rect 353 33 375 36
rect 329 28 332 33
rect 354 28 357 33
rect 368 32 374 33
rect 383 28 386 43
rect 390 36 393 37
rect 389 33 396 36
rect 404 36 407 43
rect 404 33 412 36
rect 420 36 423 43
rect 427 36 430 43
rect 420 33 430 36
rect 389 32 395 33
rect 404 28 407 33
rect 420 28 423 33
rect 427 28 430 33
rect 436 38 439 43
rect 436 37 441 38
rect 436 34 447 37
rect 455 36 458 44
rect 462 51 465 61
rect 480 54 487 58
rect 507 54 508 58
rect 522 52 525 61
rect 480 37 483 43
rect 436 28 439 34
rect 455 33 463 36
rect 479 36 483 37
rect 497 36 500 43
rect 479 33 500 36
rect 455 28 458 33
rect 480 28 483 33
rect 497 28 500 33
rect 506 37 509 43
rect 515 37 519 38
rect 506 34 523 37
rect 531 36 534 44
rect 538 51 541 61
rect 556 54 562 58
rect 576 51 579 61
rect 597 51 600 61
rect 613 51 616 61
rect 639 54 640 58
rect 648 52 651 61
rect 556 37 559 43
rect 506 28 509 34
rect 531 33 539 36
rect 555 36 559 37
rect 571 36 574 37
rect 555 33 577 36
rect 531 28 534 33
rect 556 28 559 33
rect 570 32 576 33
rect 585 28 588 43
rect 592 36 595 37
rect 591 33 598 36
rect 606 36 609 43
rect 606 33 614 36
rect 622 36 625 43
rect 629 36 632 43
rect 622 33 632 36
rect 591 32 597 33
rect 606 28 609 33
rect 622 28 625 33
rect 629 28 632 33
rect 638 38 641 43
rect 638 37 643 38
rect 638 34 649 37
rect 657 36 660 44
rect 664 51 667 61
rect 682 54 689 58
rect 709 54 710 58
rect 724 52 727 61
rect 682 37 685 43
rect 638 28 641 34
rect 657 33 665 36
rect 681 36 685 37
rect 699 36 702 43
rect 681 33 702 36
rect 657 28 660 33
rect 682 28 685 33
rect 699 28 702 33
rect 708 37 711 43
rect 717 37 721 38
rect 708 34 725 37
rect 733 36 736 44
rect 740 51 743 61
rect 758 54 764 58
rect 778 51 781 61
rect 799 51 802 61
rect 758 37 761 43
rect 708 28 711 34
rect 733 33 741 36
rect 757 36 761 37
rect 773 36 776 37
rect 757 33 779 36
rect 733 28 736 33
rect 758 28 761 33
rect 772 32 778 33
rect 787 28 790 43
rect 794 36 797 37
rect 793 33 800 36
rect 808 36 811 43
rect 808 33 818 36
rect 793 32 799 33
rect 808 28 811 33
rect 7 12 10 24
rect 24 16 25 20
rect 42 12 45 24
rect 58 12 61 24
rect 68 15 69 19
rect 94 16 95 20
rect 118 12 121 24
rect 134 12 137 24
rect 144 15 145 19
rect 172 12 175 24
rect 193 12 196 24
rect 209 12 212 24
rect 226 16 227 20
rect 244 12 247 24
rect 260 12 263 24
rect 270 15 271 19
rect 296 16 297 20
rect 320 12 323 24
rect 336 12 339 24
rect 346 15 347 19
rect 374 12 377 24
rect 395 12 398 24
rect 411 12 414 24
rect 428 16 429 20
rect 446 12 449 24
rect 462 12 465 24
rect 472 15 473 19
rect 498 16 499 20
rect 522 12 525 24
rect 538 12 541 24
rect 548 15 549 19
rect 576 12 579 24
rect 597 12 600 24
rect 613 12 616 24
rect 630 16 631 20
rect 648 12 651 24
rect 664 12 667 24
rect 674 15 675 19
rect 700 16 701 20
rect 724 12 727 24
rect 740 12 743 24
rect 750 15 751 19
rect 778 12 781 24
rect 799 12 802 24
rect 4 8 18 12
rect 22 8 38 12
rect 42 8 51 12
rect 55 8 88 12
rect 92 8 110 12
rect 114 8 127 12
rect 131 8 162 12
rect 166 8 205 12
rect 209 8 220 12
rect 224 8 240 12
rect 244 8 253 12
rect 257 8 290 12
rect 294 8 312 12
rect 316 8 329 12
rect 333 8 364 12
rect 368 8 407 12
rect 411 8 422 12
rect 426 8 442 12
rect 446 8 455 12
rect 459 8 492 12
rect 496 8 514 12
rect 518 8 531 12
rect 535 8 566 12
rect 570 8 609 12
rect 613 8 624 12
rect 628 8 644 12
rect 648 8 657 12
rect 661 8 694 12
rect 698 8 716 12
rect 720 8 733 12
rect 737 8 768 12
rect 772 8 811 12
rect 0 0 20 4
rect 24 0 84 4
rect 88 0 105 4
rect 109 0 159 4
rect 163 0 222 4
rect 226 0 286 4
rect 290 0 307 4
rect 311 0 361 4
rect 365 0 424 4
rect 428 0 488 4
rect 492 0 509 4
rect 513 0 563 4
rect 567 0 626 4
rect 630 0 690 4
rect 694 0 711 4
rect 715 0 765 4
rect 769 0 811 4
<< m2contact >>
rect 34 70 38 74
rect 61 70 65 74
rect 90 70 94 74
rect 137 70 141 74
rect 236 70 240 74
rect 263 70 267 74
rect 292 70 296 74
rect 339 70 343 74
rect 438 70 442 74
rect 465 70 469 74
rect 494 70 498 74
rect 541 70 545 74
rect 640 70 644 74
rect 667 70 671 74
rect 696 70 700 74
rect 743 70 747 74
rect 34 54 38 58
rect 83 54 87 58
rect 104 54 108 58
rect 158 54 162 58
rect 236 54 240 58
rect 285 54 289 58
rect 306 54 310 58
rect 360 54 364 58
rect 438 54 442 58
rect 487 54 491 58
rect 508 54 512 58
rect 562 54 566 58
rect 640 54 644 58
rect 689 54 693 58
rect 710 54 714 58
rect 764 54 768 58
rect 20 16 24 20
rect 64 15 68 19
rect 90 16 94 20
rect 140 15 144 19
rect 222 16 226 20
rect 266 15 270 19
rect 292 16 296 20
rect 342 15 346 19
rect 424 16 428 20
rect 468 15 472 19
rect 494 16 498 20
rect 544 15 548 19
rect 626 16 630 20
rect 670 15 674 19
rect 696 16 700 20
rect 746 15 750 19
rect 20 0 24 4
rect 84 0 88 4
rect 105 0 109 4
rect 159 0 163 4
rect 222 0 226 4
rect 286 0 290 4
rect 307 0 311 4
rect 361 0 365 4
rect 424 0 428 4
rect 488 0 492 4
rect 509 0 513 4
rect 563 0 567 4
rect 626 0 630 4
rect 690 0 694 4
rect 711 0 715 4
rect 765 0 769 4
<< metal2 >>
rect 34 58 38 70
rect 38 34 39 37
rect 20 4 24 16
rect 61 15 64 70
rect 84 4 87 54
rect 90 20 93 70
rect 105 4 108 54
rect 137 15 140 70
rect 236 58 240 70
rect 159 4 162 54
rect 165 33 166 36
rect 240 34 241 37
rect 222 4 226 16
rect 263 15 266 70
rect 286 4 289 54
rect 292 20 295 70
rect 307 4 310 54
rect 339 15 342 70
rect 438 58 442 70
rect 361 4 364 54
rect 367 33 368 36
rect 442 34 443 37
rect 424 4 428 16
rect 465 15 468 70
rect 488 4 491 54
rect 494 20 497 70
rect 509 4 512 54
rect 541 15 544 70
rect 640 58 644 70
rect 563 4 566 54
rect 569 33 570 36
rect 644 34 645 37
rect 626 4 630 16
rect 667 15 670 70
rect 690 4 693 54
rect 696 20 699 70
rect 711 4 714 54
rect 743 15 746 70
rect 765 4 768 54
rect 771 33 772 36
<< m3contact >>
rect 33 34 38 39
rect 75 33 80 38
rect 111 34 116 39
rect 151 33 156 38
rect 166 32 171 37
rect 187 32 192 37
rect 235 34 240 39
rect 277 33 282 38
rect 313 34 318 39
rect 353 33 358 38
rect 368 32 373 37
rect 389 32 394 37
rect 437 34 442 39
rect 479 33 484 38
rect 515 34 520 39
rect 555 33 560 38
rect 570 32 575 37
rect 591 32 596 37
rect 639 34 644 39
rect 681 33 686 38
rect 717 34 722 39
rect 757 33 762 38
rect 772 32 777 37
rect 793 32 798 37
<< metal3 >>
rect 111 43 192 48
rect 111 40 116 43
rect 32 39 39 40
rect 110 39 117 40
rect 32 34 33 39
rect 38 38 81 39
rect 38 34 75 38
rect 32 33 39 34
rect 74 33 75 34
rect 80 33 81 38
rect 110 34 111 39
rect 116 38 157 39
rect 187 38 192 43
rect 313 43 394 48
rect 313 40 318 43
rect 234 39 241 40
rect 312 39 319 40
rect 116 34 151 38
rect 110 33 117 34
rect 150 33 151 34
rect 156 33 157 38
rect 74 32 81 33
rect 111 27 116 33
rect 150 32 157 33
rect 165 37 172 38
rect 165 32 166 37
rect 171 32 172 37
rect 165 31 172 32
rect 186 37 193 38
rect 186 32 187 37
rect 192 32 193 37
rect 234 34 235 39
rect 240 38 283 39
rect 240 34 277 38
rect 234 33 241 34
rect 276 33 277 34
rect 282 33 283 38
rect 312 34 313 39
rect 318 38 359 39
rect 389 38 394 43
rect 515 43 596 48
rect 515 40 520 43
rect 436 39 443 40
rect 514 39 521 40
rect 318 34 353 38
rect 312 33 319 34
rect 352 33 353 34
rect 358 33 359 38
rect 276 32 283 33
rect 186 31 193 32
rect 166 27 171 31
rect 111 22 171 27
rect 313 27 318 33
rect 352 32 359 33
rect 367 37 374 38
rect 367 32 368 37
rect 373 32 374 37
rect 367 31 374 32
rect 388 37 395 38
rect 388 32 389 37
rect 394 32 395 37
rect 436 34 437 39
rect 442 38 485 39
rect 442 34 479 38
rect 436 33 443 34
rect 478 33 479 34
rect 484 33 485 38
rect 514 34 515 39
rect 520 38 561 39
rect 591 38 596 43
rect 717 43 798 48
rect 717 40 722 43
rect 638 39 645 40
rect 716 39 723 40
rect 520 34 555 38
rect 514 33 521 34
rect 554 33 555 34
rect 560 33 561 38
rect 478 32 485 33
rect 388 31 395 32
rect 368 27 373 31
rect 313 22 373 27
rect 515 27 520 33
rect 554 32 561 33
rect 569 37 576 38
rect 569 32 570 37
rect 575 32 576 37
rect 569 31 576 32
rect 590 37 597 38
rect 590 32 591 37
rect 596 32 597 37
rect 638 34 639 39
rect 644 38 687 39
rect 644 34 681 38
rect 638 33 645 34
rect 680 33 681 34
rect 686 33 687 38
rect 716 34 717 39
rect 722 38 763 39
rect 793 38 798 43
rect 722 34 757 38
rect 716 33 723 34
rect 756 33 757 34
rect 762 33 763 38
rect 680 32 687 33
rect 590 31 597 32
rect 570 27 575 31
rect 515 22 575 27
rect 717 27 722 33
rect 756 32 763 33
rect 771 37 778 38
rect 771 32 772 37
rect 777 32 778 37
rect 771 31 778 32
rect 792 37 799 38
rect 792 32 793 37
rect 798 32 799 37
rect 792 31 799 32
rect 772 27 777 31
rect 717 22 777 27
<< labels >>
rlabel metal1 3 33 7 36 1 D
rlabel metal1 181 31 184 38 1 ~Q0
rlabel metal1 202 31 205 38 1 Q0
rlabel metal1 383 31 386 38 1 ~Q1
rlabel metal1 404 31 407 38 1 Q1
rlabel metal1 0 70 10 74 4 phi
rlabel metal1 0 0 10 4 2 ~phi
rlabel metal1 4 8 14 12 1 GND!
rlabel metal1 5 61 15 65 1 Vdd!
rlabel metal1 407 70 417 74 4 phi
rlabel metal1 407 0 417 4 2 ~phi
rlabel metal1 411 8 421 12 1 GND!
rlabel metal1 412 61 422 65 1 Vdd!
rlabel metal1 585 31 588 38 1 ~Q2
rlabel metal1 606 31 609 38 1 Q2
rlabel metal1 787 31 790 38 1 ~Q3
rlabel metal1 808 31 811 38 1 Q3
<< end >>
