magic
tech scmos
timestamp 1608104093
<< ntransistor >>
rect 101 191 103 195
rect 106 191 108 195
rect 122 191 124 195
rect 138 191 140 195
rect 143 191 145 195
rect 164 191 166 195
rect 180 191 182 195
rect 196 191 198 195
rect 201 191 203 195
rect 217 191 219 195
rect 233 191 235 195
rect 238 191 240 195
rect 254 191 256 195
rect 270 191 272 195
rect 275 191 277 195
rect 296 191 298 195
rect 312 191 314 195
rect 328 191 330 195
rect 333 191 335 195
rect 349 191 351 195
rect 365 191 367 195
rect 370 191 372 195
rect 386 191 388 195
rect 402 191 404 195
rect 407 191 409 195
rect 428 191 430 195
rect 444 191 446 195
rect 460 191 462 195
rect 465 191 467 195
rect 481 191 483 195
rect 216 147 218 151
rect 240 147 242 151
rect 236 136 238 140
rect 227 122 231 124
rect 216 113 218 117
rect 240 113 242 117
rect 101 51 103 55
rect 106 51 108 55
rect 122 51 124 55
rect 138 51 140 55
rect 143 51 145 55
rect 164 51 166 55
rect 180 51 182 55
rect 196 51 198 55
rect 201 51 203 55
rect 217 51 219 55
rect 233 51 235 55
rect 238 51 240 55
rect 254 51 256 55
rect 270 51 272 55
rect 275 51 277 55
rect 296 51 298 55
rect 312 51 314 55
rect 328 51 330 55
rect 333 51 335 55
rect 349 51 351 55
rect 365 51 367 55
rect 370 51 372 55
rect 386 51 388 55
rect 402 51 404 55
rect 407 51 409 55
rect 428 51 430 55
rect 444 51 446 55
rect 460 51 462 55
rect 465 51 467 55
rect 481 51 483 55
rect 101 -35 103 -31
rect 106 -35 108 -31
rect 122 -35 124 -31
rect 138 -35 140 -31
rect 143 -35 145 -31
rect 164 -35 166 -31
rect 180 -35 182 -31
rect 196 -35 198 -31
rect 201 -35 203 -31
rect 217 -35 219 -31
rect 233 -35 235 -31
rect 238 -35 240 -31
rect 254 -35 256 -31
rect 270 -35 272 -31
rect 275 -35 277 -31
rect 296 -35 298 -31
rect 312 -35 314 -31
rect 328 -35 330 -31
rect 333 -35 335 -31
rect 349 -35 351 -31
rect 365 -35 367 -31
rect 370 -35 372 -31
rect 386 -35 388 -31
rect 402 -35 404 -31
rect 407 -35 409 -31
rect 428 -35 430 -31
rect 444 -35 446 -31
rect 460 -35 462 -31
rect 465 -35 467 -31
rect 481 -35 483 -31
rect 333 -79 335 -75
rect 357 -79 359 -75
rect 353 -90 355 -86
rect 344 -104 348 -102
rect 333 -113 335 -109
rect 357 -113 359 -109
rect 101 -175 103 -171
rect 106 -175 108 -171
rect 122 -175 124 -171
rect 138 -175 140 -171
rect 143 -175 145 -171
rect 164 -175 166 -171
rect 180 -175 182 -171
rect 196 -175 198 -171
rect 201 -175 203 -171
rect 217 -175 219 -171
rect 233 -175 235 -171
rect 238 -175 240 -171
rect 254 -175 256 -171
rect 270 -175 272 -171
rect 275 -175 277 -171
rect 296 -175 298 -171
rect 312 -175 314 -171
rect 328 -175 330 -171
rect 333 -175 335 -171
rect 349 -175 351 -171
rect 365 -175 367 -171
rect 370 -175 372 -171
rect 386 -175 388 -171
rect 402 -175 404 -171
rect 407 -175 409 -171
rect 428 -175 430 -171
rect 444 -175 446 -171
rect 460 -175 462 -171
rect 465 -175 467 -171
rect 481 -175 483 -171
<< ptransistor >>
rect 101 214 103 222
rect 106 214 108 222
rect 122 214 124 222
rect 138 214 140 222
rect 143 214 145 222
rect 164 214 166 222
rect 180 214 182 222
rect 196 214 198 222
rect 201 214 203 222
rect 217 214 219 222
rect 233 214 235 222
rect 238 214 240 222
rect 254 214 256 222
rect 270 214 272 222
rect 275 214 277 222
rect 296 214 298 222
rect 312 214 314 222
rect 328 214 330 222
rect 333 214 335 222
rect 349 214 351 222
rect 365 214 367 222
rect 370 214 372 222
rect 386 214 388 222
rect 402 214 404 222
rect 407 214 409 222
rect 428 214 430 222
rect 444 214 446 222
rect 460 214 462 222
rect 465 214 467 222
rect 481 214 483 222
rect 101 74 103 82
rect 106 74 108 82
rect 122 74 124 82
rect 138 74 140 82
rect 143 74 145 82
rect 164 74 166 82
rect 180 74 182 82
rect 196 74 198 82
rect 201 74 203 82
rect 217 74 219 82
rect 233 74 235 82
rect 238 74 240 82
rect 254 74 256 82
rect 270 74 272 82
rect 275 74 277 82
rect 296 74 298 82
rect 312 74 314 82
rect 328 74 330 82
rect 333 74 335 82
rect 349 74 351 82
rect 365 74 367 82
rect 370 74 372 82
rect 386 74 388 82
rect 402 74 404 82
rect 407 74 409 82
rect 428 74 430 82
rect 444 74 446 82
rect 460 74 462 82
rect 465 74 467 82
rect 481 74 483 82
rect 101 -12 103 -4
rect 106 -12 108 -4
rect 122 -12 124 -4
rect 138 -12 140 -4
rect 143 -12 145 -4
rect 164 -12 166 -4
rect 180 -12 182 -4
rect 196 -12 198 -4
rect 201 -12 203 -4
rect 217 -12 219 -4
rect 233 -12 235 -4
rect 238 -12 240 -4
rect 254 -12 256 -4
rect 270 -12 272 -4
rect 275 -12 277 -4
rect 296 -12 298 -4
rect 312 -12 314 -4
rect 328 -12 330 -4
rect 333 -12 335 -4
rect 349 -12 351 -4
rect 365 -12 367 -4
rect 370 -12 372 -4
rect 386 -12 388 -4
rect 402 -12 404 -4
rect 407 -12 409 -4
rect 428 -12 430 -4
rect 444 -12 446 -4
rect 460 -12 462 -4
rect 465 -12 467 -4
rect 481 -12 483 -4
rect 101 -152 103 -144
rect 106 -152 108 -144
rect 122 -152 124 -144
rect 138 -152 140 -144
rect 143 -152 145 -144
rect 164 -152 166 -144
rect 180 -152 182 -144
rect 196 -152 198 -144
rect 201 -152 203 -144
rect 217 -152 219 -144
rect 233 -152 235 -144
rect 238 -152 240 -144
rect 254 -152 256 -144
rect 270 -152 272 -144
rect 275 -152 277 -144
rect 296 -152 298 -144
rect 312 -152 314 -144
rect 328 -152 330 -144
rect 333 -152 335 -144
rect 349 -152 351 -144
rect 365 -152 367 -144
rect 370 -152 372 -144
rect 386 -152 388 -144
rect 402 -152 404 -144
rect 407 -152 409 -144
rect 428 -152 430 -144
rect 444 -152 446 -144
rect 460 -152 462 -144
rect 465 -152 467 -144
rect 481 -152 483 -144
<< ndiffusion >>
rect 100 191 101 195
rect 103 191 106 195
rect 108 191 109 195
rect 121 191 122 195
rect 124 191 125 195
rect 137 191 138 195
rect 140 191 143 195
rect 145 191 146 195
rect 163 191 164 195
rect 166 191 167 195
rect 179 191 180 195
rect 182 191 183 195
rect 195 191 196 195
rect 198 191 201 195
rect 203 191 204 195
rect 216 191 217 195
rect 219 191 220 195
rect 232 191 233 195
rect 235 191 238 195
rect 240 191 241 195
rect 253 191 254 195
rect 256 191 257 195
rect 269 191 270 195
rect 272 191 275 195
rect 277 191 278 195
rect 295 191 296 195
rect 298 191 299 195
rect 311 191 312 195
rect 314 191 315 195
rect 327 191 328 195
rect 330 191 333 195
rect 335 191 336 195
rect 348 191 349 195
rect 351 191 352 195
rect 364 191 365 195
rect 367 191 370 195
rect 372 191 373 195
rect 385 191 386 195
rect 388 191 389 195
rect 401 191 402 195
rect 404 191 407 195
rect 409 191 410 195
rect 427 191 428 195
rect 430 191 431 195
rect 443 191 444 195
rect 446 191 447 195
rect 459 191 460 195
rect 462 191 465 195
rect 467 191 468 195
rect 480 191 481 195
rect 483 191 484 195
rect 215 147 216 151
rect 218 147 219 151
rect 239 147 240 151
rect 242 147 243 151
rect 235 136 236 140
rect 238 136 239 140
rect 227 124 231 125
rect 227 121 231 122
rect 215 113 216 117
rect 218 113 219 117
rect 239 113 240 117
rect 242 113 243 117
rect 100 51 101 55
rect 103 51 106 55
rect 108 51 109 55
rect 121 51 122 55
rect 124 51 125 55
rect 137 51 138 55
rect 140 51 143 55
rect 145 51 146 55
rect 163 51 164 55
rect 166 51 167 55
rect 179 51 180 55
rect 182 51 183 55
rect 195 51 196 55
rect 198 51 201 55
rect 203 51 204 55
rect 216 51 217 55
rect 219 51 220 55
rect 232 51 233 55
rect 235 51 238 55
rect 240 51 241 55
rect 253 51 254 55
rect 256 51 257 55
rect 269 51 270 55
rect 272 51 275 55
rect 277 51 278 55
rect 295 51 296 55
rect 298 51 299 55
rect 311 51 312 55
rect 314 51 315 55
rect 327 51 328 55
rect 330 51 333 55
rect 335 51 336 55
rect 348 51 349 55
rect 351 51 352 55
rect 364 51 365 55
rect 367 51 370 55
rect 372 51 373 55
rect 385 51 386 55
rect 388 51 389 55
rect 401 51 402 55
rect 404 51 407 55
rect 409 51 410 55
rect 427 51 428 55
rect 430 51 431 55
rect 443 51 444 55
rect 446 51 447 55
rect 459 51 460 55
rect 462 51 465 55
rect 467 51 468 55
rect 480 51 481 55
rect 483 51 484 55
rect 100 -35 101 -31
rect 103 -35 106 -31
rect 108 -35 109 -31
rect 121 -35 122 -31
rect 124 -35 125 -31
rect 137 -35 138 -31
rect 140 -35 143 -31
rect 145 -35 146 -31
rect 163 -35 164 -31
rect 166 -35 167 -31
rect 179 -35 180 -31
rect 182 -35 183 -31
rect 195 -35 196 -31
rect 198 -35 201 -31
rect 203 -35 204 -31
rect 216 -35 217 -31
rect 219 -35 220 -31
rect 232 -35 233 -31
rect 235 -35 238 -31
rect 240 -35 241 -31
rect 253 -35 254 -31
rect 256 -35 257 -31
rect 269 -35 270 -31
rect 272 -35 275 -31
rect 277 -35 278 -31
rect 295 -35 296 -31
rect 298 -35 299 -31
rect 311 -35 312 -31
rect 314 -35 315 -31
rect 327 -35 328 -31
rect 330 -35 333 -31
rect 335 -35 336 -31
rect 348 -35 349 -31
rect 351 -35 352 -31
rect 364 -35 365 -31
rect 367 -35 370 -31
rect 372 -35 373 -31
rect 385 -35 386 -31
rect 388 -35 389 -31
rect 401 -35 402 -31
rect 404 -35 407 -31
rect 409 -35 410 -31
rect 427 -35 428 -31
rect 430 -35 431 -31
rect 443 -35 444 -31
rect 446 -35 447 -31
rect 459 -35 460 -31
rect 462 -35 465 -31
rect 467 -35 468 -31
rect 480 -35 481 -31
rect 483 -35 484 -31
rect 332 -79 333 -75
rect 335 -79 336 -75
rect 356 -79 357 -75
rect 359 -79 360 -75
rect 352 -90 353 -86
rect 355 -90 356 -86
rect 344 -102 348 -101
rect 344 -105 348 -104
rect 332 -113 333 -109
rect 335 -113 336 -109
rect 356 -113 357 -109
rect 359 -113 360 -109
rect 100 -175 101 -171
rect 103 -175 106 -171
rect 108 -175 109 -171
rect 121 -175 122 -171
rect 124 -175 125 -171
rect 137 -175 138 -171
rect 140 -175 143 -171
rect 145 -175 146 -171
rect 163 -175 164 -171
rect 166 -175 167 -171
rect 179 -175 180 -171
rect 182 -175 183 -171
rect 195 -175 196 -171
rect 198 -175 201 -171
rect 203 -175 204 -171
rect 216 -175 217 -171
rect 219 -175 220 -171
rect 232 -175 233 -171
rect 235 -175 238 -171
rect 240 -175 241 -171
rect 253 -175 254 -171
rect 256 -175 257 -171
rect 269 -175 270 -171
rect 272 -175 275 -171
rect 277 -175 278 -171
rect 295 -175 296 -171
rect 298 -175 299 -171
rect 311 -175 312 -171
rect 314 -175 315 -171
rect 327 -175 328 -171
rect 330 -175 333 -171
rect 335 -175 336 -171
rect 348 -175 349 -171
rect 351 -175 352 -171
rect 364 -175 365 -171
rect 367 -175 370 -171
rect 372 -175 373 -171
rect 385 -175 386 -171
rect 388 -175 389 -171
rect 401 -175 402 -171
rect 404 -175 407 -171
rect 409 -175 410 -171
rect 427 -175 428 -171
rect 430 -175 431 -171
rect 443 -175 444 -171
rect 446 -175 447 -171
rect 459 -175 460 -171
rect 462 -175 465 -171
rect 467 -175 468 -171
rect 480 -175 481 -171
rect 483 -175 484 -171
<< pdiffusion >>
rect 100 214 101 222
rect 103 214 106 222
rect 108 214 109 222
rect 121 214 122 222
rect 124 218 125 222
rect 124 214 129 218
rect 137 214 138 222
rect 140 214 143 222
rect 145 214 146 222
rect 163 214 164 222
rect 166 214 167 222
rect 179 214 180 222
rect 182 218 183 222
rect 182 214 187 218
rect 195 214 196 222
rect 198 214 201 222
rect 203 214 204 222
rect 216 214 217 222
rect 219 214 220 222
rect 232 214 233 222
rect 235 214 238 222
rect 240 214 241 222
rect 253 214 254 222
rect 256 218 257 222
rect 256 214 261 218
rect 269 214 270 222
rect 272 214 275 222
rect 277 214 278 222
rect 295 214 296 222
rect 298 214 299 222
rect 311 214 312 222
rect 314 218 315 222
rect 314 214 319 218
rect 327 214 328 222
rect 330 214 333 222
rect 335 214 336 222
rect 348 214 349 222
rect 351 214 352 222
rect 364 214 365 222
rect 367 214 370 222
rect 372 214 373 222
rect 385 214 386 222
rect 388 218 389 222
rect 388 214 393 218
rect 401 214 402 222
rect 404 214 407 222
rect 409 214 410 222
rect 427 214 428 222
rect 430 214 431 222
rect 443 214 444 222
rect 446 218 447 222
rect 446 214 451 218
rect 459 214 460 222
rect 462 214 465 222
rect 467 214 468 222
rect 480 214 481 222
rect 483 214 484 222
rect 100 74 101 82
rect 103 74 106 82
rect 108 74 109 82
rect 121 74 122 82
rect 124 78 125 82
rect 124 74 129 78
rect 137 74 138 82
rect 140 74 143 82
rect 145 74 146 82
rect 163 74 164 82
rect 166 74 167 82
rect 179 74 180 82
rect 182 78 183 82
rect 182 74 187 78
rect 195 74 196 82
rect 198 74 201 82
rect 203 74 204 82
rect 216 74 217 82
rect 219 74 220 82
rect 232 74 233 82
rect 235 74 238 82
rect 240 74 241 82
rect 253 74 254 82
rect 256 78 257 82
rect 256 74 261 78
rect 269 74 270 82
rect 272 74 275 82
rect 277 74 278 82
rect 295 74 296 82
rect 298 74 299 82
rect 311 74 312 82
rect 314 78 315 82
rect 314 74 319 78
rect 327 74 328 82
rect 330 74 333 82
rect 335 74 336 82
rect 348 74 349 82
rect 351 74 352 82
rect 364 74 365 82
rect 367 74 370 82
rect 372 74 373 82
rect 385 74 386 82
rect 388 78 389 82
rect 388 74 393 78
rect 401 74 402 82
rect 404 74 407 82
rect 409 74 410 82
rect 427 74 428 82
rect 430 74 431 82
rect 443 74 444 82
rect 446 78 447 82
rect 446 74 451 78
rect 459 74 460 82
rect 462 74 465 82
rect 467 74 468 82
rect 480 74 481 82
rect 483 74 484 82
rect 100 -12 101 -4
rect 103 -12 106 -4
rect 108 -12 109 -4
rect 121 -12 122 -4
rect 124 -8 125 -4
rect 124 -12 129 -8
rect 137 -12 138 -4
rect 140 -12 143 -4
rect 145 -12 146 -4
rect 163 -12 164 -4
rect 166 -12 167 -4
rect 179 -12 180 -4
rect 182 -8 183 -4
rect 182 -12 187 -8
rect 195 -12 196 -4
rect 198 -12 201 -4
rect 203 -12 204 -4
rect 216 -12 217 -4
rect 219 -12 220 -4
rect 232 -12 233 -4
rect 235 -12 238 -4
rect 240 -12 241 -4
rect 253 -12 254 -4
rect 256 -8 257 -4
rect 256 -12 261 -8
rect 269 -12 270 -4
rect 272 -12 275 -4
rect 277 -12 278 -4
rect 295 -12 296 -4
rect 298 -12 299 -4
rect 311 -12 312 -4
rect 314 -8 315 -4
rect 314 -12 319 -8
rect 327 -12 328 -4
rect 330 -12 333 -4
rect 335 -12 336 -4
rect 348 -12 349 -4
rect 351 -12 352 -4
rect 364 -12 365 -4
rect 367 -12 370 -4
rect 372 -12 373 -4
rect 385 -12 386 -4
rect 388 -8 389 -4
rect 388 -12 393 -8
rect 401 -12 402 -4
rect 404 -12 407 -4
rect 409 -12 410 -4
rect 427 -12 428 -4
rect 430 -12 431 -4
rect 443 -12 444 -4
rect 446 -8 447 -4
rect 446 -12 451 -8
rect 459 -12 460 -4
rect 462 -12 465 -4
rect 467 -12 468 -4
rect 480 -12 481 -4
rect 483 -12 484 -4
rect 100 -152 101 -144
rect 103 -152 106 -144
rect 108 -152 109 -144
rect 121 -152 122 -144
rect 124 -148 125 -144
rect 124 -152 129 -148
rect 137 -152 138 -144
rect 140 -152 143 -144
rect 145 -152 146 -144
rect 163 -152 164 -144
rect 166 -152 167 -144
rect 179 -152 180 -144
rect 182 -148 183 -144
rect 182 -152 187 -148
rect 195 -152 196 -144
rect 198 -152 201 -144
rect 203 -152 204 -144
rect 216 -152 217 -144
rect 219 -152 220 -144
rect 232 -152 233 -144
rect 235 -152 238 -144
rect 240 -152 241 -144
rect 253 -152 254 -144
rect 256 -148 257 -144
rect 256 -152 261 -148
rect 269 -152 270 -144
rect 272 -152 275 -144
rect 277 -152 278 -144
rect 295 -152 296 -144
rect 298 -152 299 -144
rect 311 -152 312 -144
rect 314 -148 315 -144
rect 314 -152 319 -148
rect 327 -152 328 -144
rect 330 -152 333 -144
rect 335 -152 336 -144
rect 348 -152 349 -144
rect 351 -152 352 -144
rect 364 -152 365 -144
rect 367 -152 370 -144
rect 372 -152 373 -144
rect 385 -152 386 -144
rect 388 -148 389 -144
rect 388 -152 393 -148
rect 401 -152 402 -144
rect 404 -152 407 -144
rect 409 -152 410 -144
rect 427 -152 428 -144
rect 430 -152 431 -144
rect 443 -152 444 -144
rect 446 -148 447 -144
rect 446 -152 451 -148
rect 459 -152 460 -144
rect 462 -152 465 -144
rect 467 -152 468 -144
rect 480 -152 481 -144
rect 483 -152 484 -144
<< ndcontact >>
rect 96 191 100 195
rect 109 191 113 195
rect 117 191 121 195
rect 125 191 129 195
rect 133 191 137 195
rect 146 191 150 195
rect 159 191 163 195
rect 167 191 171 195
rect 175 191 179 195
rect 183 191 187 195
rect 191 191 195 195
rect 204 191 208 195
rect 212 191 216 195
rect 220 191 224 195
rect 228 191 232 195
rect 241 191 245 195
rect 249 191 253 195
rect 257 191 261 195
rect 265 191 269 195
rect 278 191 282 195
rect 291 191 295 195
rect 299 191 303 195
rect 307 191 311 195
rect 315 191 319 195
rect 323 191 327 195
rect 336 191 340 195
rect 344 191 348 195
rect 352 191 356 195
rect 360 191 364 195
rect 373 191 377 195
rect 381 191 385 195
rect 389 191 393 195
rect 397 191 401 195
rect 410 191 414 195
rect 423 191 427 195
rect 431 191 435 195
rect 439 191 443 195
rect 447 191 451 195
rect 455 191 459 195
rect 468 191 472 195
rect 476 191 480 195
rect 484 191 488 195
rect 211 147 215 151
rect 219 147 223 151
rect 235 147 239 151
rect 243 147 247 151
rect 231 136 235 140
rect 239 136 243 140
rect 227 125 231 129
rect 227 117 231 121
rect 211 113 215 117
rect 219 113 223 117
rect 235 113 239 117
rect 243 113 247 117
rect 96 51 100 55
rect 109 51 113 55
rect 117 51 121 55
rect 125 51 129 55
rect 133 51 137 55
rect 146 51 150 55
rect 159 51 163 55
rect 167 51 171 55
rect 175 51 179 55
rect 183 51 187 55
rect 191 51 195 55
rect 204 51 208 55
rect 212 51 216 55
rect 220 51 224 55
rect 228 51 232 55
rect 241 51 245 55
rect 249 51 253 55
rect 257 51 261 55
rect 265 51 269 55
rect 278 51 282 55
rect 291 51 295 55
rect 299 51 303 55
rect 307 51 311 55
rect 315 51 319 55
rect 323 51 327 55
rect 336 51 340 55
rect 344 51 348 55
rect 352 51 356 55
rect 360 51 364 55
rect 373 51 377 55
rect 381 51 385 55
rect 389 51 393 55
rect 397 51 401 55
rect 410 51 414 55
rect 423 51 427 55
rect 431 51 435 55
rect 439 51 443 55
rect 447 51 451 55
rect 455 51 459 55
rect 468 51 472 55
rect 476 51 480 55
rect 484 51 488 55
rect 96 -35 100 -31
rect 109 -35 113 -31
rect 117 -35 121 -31
rect 125 -35 129 -31
rect 133 -35 137 -31
rect 146 -35 150 -31
rect 159 -35 163 -31
rect 167 -35 171 -31
rect 175 -35 179 -31
rect 183 -35 187 -31
rect 191 -35 195 -31
rect 204 -35 208 -31
rect 212 -35 216 -31
rect 220 -35 224 -31
rect 228 -35 232 -31
rect 241 -35 245 -31
rect 249 -35 253 -31
rect 257 -35 261 -31
rect 265 -35 269 -31
rect 278 -35 282 -31
rect 291 -35 295 -31
rect 299 -35 303 -31
rect 307 -35 311 -31
rect 315 -35 319 -31
rect 323 -35 327 -31
rect 336 -35 340 -31
rect 344 -35 348 -31
rect 352 -35 356 -31
rect 360 -35 364 -31
rect 373 -35 377 -31
rect 381 -35 385 -31
rect 389 -35 393 -31
rect 397 -35 401 -31
rect 410 -35 414 -31
rect 423 -35 427 -31
rect 431 -35 435 -31
rect 439 -35 443 -31
rect 447 -35 451 -31
rect 455 -35 459 -31
rect 468 -35 472 -31
rect 476 -35 480 -31
rect 484 -35 488 -31
rect 328 -79 332 -75
rect 336 -79 340 -75
rect 352 -79 356 -75
rect 360 -79 364 -75
rect 348 -90 352 -86
rect 356 -90 360 -86
rect 344 -101 348 -97
rect 344 -109 348 -105
rect 328 -113 332 -109
rect 336 -113 340 -109
rect 352 -113 356 -109
rect 360 -113 364 -109
rect 96 -175 100 -171
rect 109 -175 113 -171
rect 117 -175 121 -171
rect 125 -175 129 -171
rect 133 -175 137 -171
rect 146 -175 150 -171
rect 159 -175 163 -171
rect 167 -175 171 -171
rect 175 -175 179 -171
rect 183 -175 187 -171
rect 191 -175 195 -171
rect 204 -175 208 -171
rect 212 -175 216 -171
rect 220 -175 224 -171
rect 228 -175 232 -171
rect 241 -175 245 -171
rect 249 -175 253 -171
rect 257 -175 261 -171
rect 265 -175 269 -171
rect 278 -175 282 -171
rect 291 -175 295 -171
rect 299 -175 303 -171
rect 307 -175 311 -171
rect 315 -175 319 -171
rect 323 -175 327 -171
rect 336 -175 340 -171
rect 344 -175 348 -171
rect 352 -175 356 -171
rect 360 -175 364 -171
rect 373 -175 377 -171
rect 381 -175 385 -171
rect 389 -175 393 -171
rect 397 -175 401 -171
rect 410 -175 414 -171
rect 423 -175 427 -171
rect 431 -175 435 -171
rect 439 -175 443 -171
rect 447 -175 451 -171
rect 455 -175 459 -171
rect 468 -175 472 -171
rect 476 -175 480 -171
rect 484 -175 488 -171
<< pdcontact >>
rect 96 214 100 222
rect 109 214 113 222
rect 117 214 121 222
rect 125 218 129 222
rect 133 214 137 222
rect 146 214 150 222
rect 159 214 163 222
rect 167 214 171 222
rect 175 214 179 222
rect 183 218 187 222
rect 191 214 195 222
rect 204 214 208 222
rect 212 214 216 222
rect 220 214 224 222
rect 228 214 232 222
rect 241 214 245 222
rect 249 214 253 222
rect 257 218 261 222
rect 265 214 269 222
rect 278 214 282 222
rect 291 214 295 222
rect 299 214 303 222
rect 307 214 311 222
rect 315 218 319 222
rect 323 214 327 222
rect 336 214 340 222
rect 344 214 348 222
rect 352 214 356 222
rect 360 214 364 222
rect 373 214 377 222
rect 381 214 385 222
rect 389 218 393 222
rect 397 214 401 222
rect 410 214 414 222
rect 423 214 427 222
rect 431 214 435 222
rect 439 214 443 222
rect 447 218 451 222
rect 455 214 459 222
rect 468 214 472 222
rect 476 214 480 222
rect 484 214 488 222
rect 96 74 100 82
rect 109 74 113 82
rect 117 74 121 82
rect 125 78 129 82
rect 133 74 137 82
rect 146 74 150 82
rect 159 74 163 82
rect 167 74 171 82
rect 175 74 179 82
rect 183 78 187 82
rect 191 74 195 82
rect 204 74 208 82
rect 212 74 216 82
rect 220 74 224 82
rect 228 74 232 82
rect 241 74 245 82
rect 249 74 253 82
rect 257 78 261 82
rect 265 74 269 82
rect 278 74 282 82
rect 291 74 295 82
rect 299 74 303 82
rect 307 74 311 82
rect 315 78 319 82
rect 323 74 327 82
rect 336 74 340 82
rect 344 74 348 82
rect 352 74 356 82
rect 360 74 364 82
rect 373 74 377 82
rect 381 74 385 82
rect 389 78 393 82
rect 397 74 401 82
rect 410 74 414 82
rect 423 74 427 82
rect 431 74 435 82
rect 439 74 443 82
rect 447 78 451 82
rect 455 74 459 82
rect 468 74 472 82
rect 476 74 480 82
rect 484 74 488 82
rect 96 -12 100 -4
rect 109 -12 113 -4
rect 117 -12 121 -4
rect 125 -8 129 -4
rect 133 -12 137 -4
rect 146 -12 150 -4
rect 159 -12 163 -4
rect 167 -12 171 -4
rect 175 -12 179 -4
rect 183 -8 187 -4
rect 191 -12 195 -4
rect 204 -12 208 -4
rect 212 -12 216 -4
rect 220 -12 224 -4
rect 228 -12 232 -4
rect 241 -12 245 -4
rect 249 -12 253 -4
rect 257 -8 261 -4
rect 265 -12 269 -4
rect 278 -12 282 -4
rect 291 -12 295 -4
rect 299 -12 303 -4
rect 307 -12 311 -4
rect 315 -8 319 -4
rect 323 -12 327 -4
rect 336 -12 340 -4
rect 344 -12 348 -4
rect 352 -12 356 -4
rect 360 -12 364 -4
rect 373 -12 377 -4
rect 381 -12 385 -4
rect 389 -8 393 -4
rect 397 -12 401 -4
rect 410 -12 414 -4
rect 423 -12 427 -4
rect 431 -12 435 -4
rect 439 -12 443 -4
rect 447 -8 451 -4
rect 455 -12 459 -4
rect 468 -12 472 -4
rect 476 -12 480 -4
rect 484 -12 488 -4
rect 96 -152 100 -144
rect 109 -152 113 -144
rect 117 -152 121 -144
rect 125 -148 129 -144
rect 133 -152 137 -144
rect 146 -152 150 -144
rect 159 -152 163 -144
rect 167 -152 171 -144
rect 175 -152 179 -144
rect 183 -148 187 -144
rect 191 -152 195 -144
rect 204 -152 208 -144
rect 212 -152 216 -144
rect 220 -152 224 -144
rect 228 -152 232 -144
rect 241 -152 245 -144
rect 249 -152 253 -144
rect 257 -148 261 -144
rect 265 -152 269 -144
rect 278 -152 282 -144
rect 291 -152 295 -144
rect 299 -152 303 -144
rect 307 -152 311 -144
rect 315 -148 319 -144
rect 323 -152 327 -144
rect 336 -152 340 -144
rect 344 -152 348 -144
rect 352 -152 356 -144
rect 360 -152 364 -144
rect 373 -152 377 -144
rect 381 -152 385 -144
rect 389 -148 393 -144
rect 397 -152 401 -144
rect 410 -152 414 -144
rect 423 -152 427 -144
rect 431 -152 435 -144
rect 439 -152 443 -144
rect 447 -148 451 -144
rect 455 -152 459 -144
rect 468 -152 472 -144
rect 476 -152 480 -144
rect 484 -152 488 -144
<< psubstratepcontact >>
rect 126 175 130 179
rect 154 175 158 179
rect 184 175 188 179
rect 258 175 262 179
rect 286 175 290 179
rect 316 175 320 179
rect 390 175 394 179
rect 418 175 422 179
rect 448 175 452 179
rect 126 35 130 39
rect 154 35 158 39
rect 184 35 188 39
rect 258 35 262 39
rect 286 35 290 39
rect 316 35 320 39
rect 390 35 394 39
rect 418 35 422 39
rect 448 35 452 39
rect 126 -51 130 -47
rect 154 -51 158 -47
rect 184 -51 188 -47
rect 258 -51 262 -47
rect 286 -51 290 -47
rect 316 -51 320 -47
rect 390 -51 394 -47
rect 418 -51 422 -47
rect 448 -51 452 -47
rect 126 -191 130 -187
rect 154 -191 158 -187
rect 184 -191 188 -187
rect 258 -191 262 -187
rect 286 -191 290 -187
rect 316 -191 320 -187
rect 390 -191 394 -187
rect 418 -191 422 -187
rect 448 -191 452 -187
<< nsubstratencontact >>
rect 126 232 130 236
rect 154 232 158 236
rect 184 232 188 236
rect 221 232 225 236
rect 258 232 262 236
rect 286 232 290 236
rect 316 232 320 236
rect 353 232 357 236
rect 390 232 394 236
rect 418 232 422 236
rect 448 232 452 236
rect 485 232 489 236
rect 126 92 130 96
rect 154 92 158 96
rect 184 92 188 96
rect 221 92 225 96
rect 258 92 262 96
rect 286 92 290 96
rect 316 92 320 96
rect 353 92 357 96
rect 390 92 394 96
rect 418 92 422 96
rect 448 92 452 96
rect 485 92 489 96
rect 126 6 130 10
rect 154 6 158 10
rect 184 6 188 10
rect 221 6 225 10
rect 258 6 262 10
rect 286 6 290 10
rect 316 6 320 10
rect 353 6 357 10
rect 390 6 394 10
rect 418 6 422 10
rect 448 6 452 10
rect 485 6 489 10
rect 126 -134 130 -130
rect 154 -134 158 -130
rect 184 -134 188 -130
rect 221 -134 225 -130
rect 258 -134 262 -130
rect 286 -134 290 -130
rect 316 -134 320 -130
rect 353 -134 357 -130
rect 390 -134 394 -130
rect 418 -134 422 -130
rect 448 -134 452 -130
rect 485 -134 489 -130
<< polysilicon >>
rect 101 222 103 224
rect 106 222 108 225
rect 122 222 124 224
rect 138 222 140 224
rect 143 222 145 225
rect 164 222 166 225
rect 180 222 182 225
rect 196 222 198 224
rect 201 222 203 225
rect 217 222 219 224
rect 233 222 235 224
rect 238 222 240 225
rect 254 222 256 224
rect 270 222 272 224
rect 275 222 277 225
rect 296 222 298 225
rect 312 222 314 225
rect 328 222 330 224
rect 333 222 335 225
rect 349 222 351 224
rect 365 222 367 224
rect 370 222 372 225
rect 386 222 388 224
rect 402 222 404 224
rect 407 222 409 225
rect 428 222 430 225
rect 444 222 446 225
rect 460 222 462 224
rect 465 222 467 225
rect 481 222 483 224
rect 101 209 103 214
rect 106 212 108 214
rect 101 195 103 205
rect 106 195 108 202
rect 122 195 124 214
rect 138 205 140 214
rect 143 212 145 214
rect 164 212 166 214
rect 180 211 182 214
rect 138 195 140 198
rect 143 195 145 197
rect 164 195 166 197
rect 180 195 182 207
rect 196 205 198 214
rect 201 212 203 214
rect 196 195 198 198
rect 201 195 203 197
rect 217 195 219 214
rect 233 211 235 214
rect 238 212 240 214
rect 233 195 235 207
rect 238 195 240 202
rect 254 195 256 214
rect 270 205 272 214
rect 275 212 277 214
rect 296 212 298 214
rect 312 211 314 214
rect 270 195 272 198
rect 275 195 277 197
rect 296 195 298 197
rect 312 195 314 207
rect 328 205 330 214
rect 333 212 335 214
rect 328 195 330 198
rect 333 195 335 197
rect 349 195 351 214
rect 365 211 367 214
rect 370 212 372 214
rect 365 195 367 207
rect 370 195 372 202
rect 386 195 388 214
rect 402 205 404 214
rect 407 212 409 214
rect 428 212 430 214
rect 444 211 446 214
rect 402 195 404 198
rect 407 195 409 197
rect 428 195 430 197
rect 444 195 446 207
rect 460 205 462 214
rect 465 212 467 214
rect 481 206 483 214
rect 460 195 462 198
rect 465 195 467 197
rect 481 195 483 202
rect 101 189 103 191
rect 106 188 108 191
rect 122 189 124 191
rect 138 189 140 191
rect 143 186 145 191
rect 164 186 166 191
rect 180 189 182 191
rect 196 189 198 191
rect 201 186 203 191
rect 217 189 219 191
rect 233 189 235 191
rect 238 188 240 191
rect 254 189 256 191
rect 270 189 272 191
rect 275 186 277 191
rect 296 186 298 191
rect 312 189 314 191
rect 328 189 330 191
rect 333 186 335 191
rect 349 189 351 191
rect 365 189 367 191
rect 370 188 372 191
rect 386 189 388 191
rect 402 189 404 191
rect 407 186 409 191
rect 428 186 430 191
rect 444 189 446 191
rect 460 189 462 191
rect 465 186 467 191
rect 481 189 483 191
rect 216 151 218 154
rect 240 151 242 154
rect 216 145 218 147
rect 240 145 242 147
rect 236 140 238 142
rect 236 133 238 136
rect 225 122 227 124
rect 231 122 250 124
rect 216 117 218 119
rect 240 117 242 119
rect 216 110 218 113
rect 240 110 242 113
rect 101 82 103 84
rect 106 82 108 85
rect 122 82 124 84
rect 138 82 140 84
rect 143 82 145 85
rect 164 82 166 85
rect 180 82 182 85
rect 196 82 198 84
rect 201 82 203 85
rect 217 82 219 84
rect 233 82 235 84
rect 238 82 240 85
rect 254 82 256 84
rect 270 82 272 84
rect 275 82 277 85
rect 296 82 298 85
rect 312 82 314 85
rect 328 82 330 84
rect 333 82 335 85
rect 349 82 351 84
rect 365 82 367 84
rect 370 82 372 85
rect 386 82 388 84
rect 402 82 404 84
rect 407 82 409 85
rect 428 82 430 85
rect 444 82 446 85
rect 460 82 462 84
rect 465 82 467 85
rect 481 82 483 84
rect 101 69 103 74
rect 106 72 108 74
rect 101 55 103 65
rect 106 55 108 62
rect 122 55 124 74
rect 138 65 140 74
rect 143 72 145 74
rect 164 72 166 74
rect 180 71 182 74
rect 138 55 140 58
rect 143 55 145 57
rect 164 55 166 57
rect 180 55 182 67
rect 196 65 198 74
rect 201 72 203 74
rect 196 55 198 58
rect 201 55 203 57
rect 217 55 219 74
rect 233 71 235 74
rect 238 72 240 74
rect 233 55 235 67
rect 238 55 240 62
rect 254 55 256 74
rect 270 65 272 74
rect 275 72 277 74
rect 296 72 298 74
rect 312 71 314 74
rect 270 55 272 58
rect 275 55 277 57
rect 296 55 298 57
rect 312 55 314 67
rect 328 65 330 74
rect 333 72 335 74
rect 328 55 330 58
rect 333 55 335 57
rect 349 55 351 74
rect 365 71 367 74
rect 370 72 372 74
rect 365 55 367 67
rect 370 55 372 62
rect 386 55 388 74
rect 402 65 404 74
rect 407 72 409 74
rect 428 72 430 74
rect 444 71 446 74
rect 402 55 404 58
rect 407 55 409 57
rect 428 55 430 57
rect 444 55 446 67
rect 460 65 462 74
rect 465 72 467 74
rect 481 66 483 74
rect 460 55 462 58
rect 465 55 467 57
rect 481 55 483 62
rect 101 49 103 51
rect 106 48 108 51
rect 122 49 124 51
rect 138 49 140 51
rect 143 46 145 51
rect 164 46 166 51
rect 180 49 182 51
rect 196 49 198 51
rect 201 46 203 51
rect 217 49 219 51
rect 233 49 235 51
rect 238 48 240 51
rect 254 49 256 51
rect 270 49 272 51
rect 275 46 277 51
rect 296 46 298 51
rect 312 49 314 51
rect 328 49 330 51
rect 333 46 335 51
rect 349 49 351 51
rect 365 49 367 51
rect 370 48 372 51
rect 386 49 388 51
rect 402 49 404 51
rect 407 46 409 51
rect 428 46 430 51
rect 444 49 446 51
rect 460 49 462 51
rect 465 46 467 51
rect 481 49 483 51
rect 101 -4 103 -2
rect 106 -4 108 -1
rect 122 -4 124 -2
rect 138 -4 140 -2
rect 143 -4 145 -1
rect 164 -4 166 -1
rect 180 -4 182 -1
rect 196 -4 198 -2
rect 201 -4 203 -1
rect 217 -4 219 -2
rect 233 -4 235 -2
rect 238 -4 240 -1
rect 254 -4 256 -2
rect 270 -4 272 -2
rect 275 -4 277 -1
rect 296 -4 298 -1
rect 312 -4 314 -1
rect 328 -4 330 -2
rect 333 -4 335 -1
rect 349 -4 351 -2
rect 365 -4 367 -2
rect 370 -4 372 -1
rect 386 -4 388 -2
rect 402 -4 404 -2
rect 407 -4 409 -1
rect 428 -4 430 -1
rect 444 -4 446 -1
rect 460 -4 462 -2
rect 465 -4 467 -1
rect 481 -4 483 -2
rect 101 -17 103 -12
rect 106 -14 108 -12
rect 101 -31 103 -21
rect 106 -31 108 -24
rect 122 -31 124 -12
rect 138 -21 140 -12
rect 143 -14 145 -12
rect 164 -14 166 -12
rect 180 -15 182 -12
rect 138 -31 140 -28
rect 143 -31 145 -29
rect 164 -31 166 -29
rect 180 -31 182 -19
rect 196 -21 198 -12
rect 201 -14 203 -12
rect 196 -31 198 -28
rect 201 -31 203 -29
rect 217 -31 219 -12
rect 233 -15 235 -12
rect 238 -14 240 -12
rect 233 -31 235 -19
rect 238 -31 240 -24
rect 254 -31 256 -12
rect 270 -21 272 -12
rect 275 -14 277 -12
rect 296 -14 298 -12
rect 312 -15 314 -12
rect 270 -31 272 -28
rect 275 -31 277 -29
rect 296 -31 298 -29
rect 312 -31 314 -19
rect 328 -21 330 -12
rect 333 -14 335 -12
rect 328 -31 330 -28
rect 333 -31 335 -29
rect 349 -31 351 -12
rect 365 -15 367 -12
rect 370 -14 372 -12
rect 365 -31 367 -19
rect 370 -31 372 -24
rect 386 -31 388 -12
rect 402 -21 404 -12
rect 407 -14 409 -12
rect 428 -14 430 -12
rect 444 -15 446 -12
rect 402 -31 404 -28
rect 407 -31 409 -29
rect 428 -31 430 -29
rect 444 -31 446 -19
rect 460 -21 462 -12
rect 465 -14 467 -12
rect 481 -20 483 -12
rect 460 -31 462 -28
rect 465 -31 467 -29
rect 481 -31 483 -24
rect 101 -37 103 -35
rect 106 -38 108 -35
rect 122 -37 124 -35
rect 138 -37 140 -35
rect 143 -40 145 -35
rect 164 -40 166 -35
rect 180 -37 182 -35
rect 196 -37 198 -35
rect 201 -40 203 -35
rect 217 -37 219 -35
rect 233 -37 235 -35
rect 238 -38 240 -35
rect 254 -37 256 -35
rect 270 -37 272 -35
rect 275 -40 277 -35
rect 296 -40 298 -35
rect 312 -37 314 -35
rect 328 -37 330 -35
rect 333 -40 335 -35
rect 349 -37 351 -35
rect 365 -37 367 -35
rect 370 -38 372 -35
rect 386 -37 388 -35
rect 402 -37 404 -35
rect 407 -40 409 -35
rect 428 -40 430 -35
rect 444 -37 446 -35
rect 460 -37 462 -35
rect 465 -40 467 -35
rect 481 -37 483 -35
rect 333 -75 335 -72
rect 357 -75 359 -72
rect 333 -81 335 -79
rect 357 -81 359 -79
rect 353 -86 355 -84
rect 353 -93 355 -90
rect 342 -104 344 -102
rect 348 -104 367 -102
rect 333 -109 335 -107
rect 357 -109 359 -107
rect 333 -116 335 -113
rect 357 -116 359 -113
rect 101 -144 103 -142
rect 106 -144 108 -141
rect 122 -144 124 -142
rect 138 -144 140 -142
rect 143 -144 145 -141
rect 164 -144 166 -141
rect 180 -144 182 -141
rect 196 -144 198 -142
rect 201 -144 203 -141
rect 217 -144 219 -142
rect 233 -144 235 -142
rect 238 -144 240 -141
rect 254 -144 256 -142
rect 270 -144 272 -142
rect 275 -144 277 -141
rect 296 -144 298 -141
rect 312 -144 314 -141
rect 328 -144 330 -142
rect 333 -144 335 -141
rect 349 -144 351 -142
rect 365 -144 367 -142
rect 370 -144 372 -141
rect 386 -144 388 -142
rect 402 -144 404 -142
rect 407 -144 409 -141
rect 428 -144 430 -141
rect 444 -144 446 -141
rect 460 -144 462 -142
rect 465 -144 467 -141
rect 481 -144 483 -142
rect 101 -157 103 -152
rect 106 -154 108 -152
rect 101 -171 103 -161
rect 106 -171 108 -164
rect 122 -171 124 -152
rect 138 -161 140 -152
rect 143 -154 145 -152
rect 164 -154 166 -152
rect 180 -155 182 -152
rect 138 -171 140 -168
rect 143 -171 145 -169
rect 164 -171 166 -169
rect 180 -171 182 -159
rect 196 -161 198 -152
rect 201 -154 203 -152
rect 196 -171 198 -168
rect 201 -171 203 -169
rect 217 -171 219 -152
rect 233 -155 235 -152
rect 238 -154 240 -152
rect 233 -171 235 -159
rect 238 -171 240 -164
rect 254 -171 256 -152
rect 270 -161 272 -152
rect 275 -154 277 -152
rect 296 -154 298 -152
rect 312 -155 314 -152
rect 270 -171 272 -168
rect 275 -171 277 -169
rect 296 -171 298 -169
rect 312 -171 314 -159
rect 328 -161 330 -152
rect 333 -154 335 -152
rect 328 -171 330 -168
rect 333 -171 335 -169
rect 349 -171 351 -152
rect 365 -155 367 -152
rect 370 -154 372 -152
rect 365 -171 367 -159
rect 370 -171 372 -164
rect 386 -171 388 -152
rect 402 -161 404 -152
rect 407 -154 409 -152
rect 428 -154 430 -152
rect 444 -155 446 -152
rect 402 -171 404 -168
rect 407 -171 409 -169
rect 428 -171 430 -169
rect 444 -171 446 -159
rect 460 -161 462 -152
rect 465 -154 467 -152
rect 481 -160 483 -152
rect 460 -171 462 -168
rect 465 -171 467 -169
rect 481 -171 483 -164
rect 101 -177 103 -175
rect 106 -178 108 -175
rect 122 -177 124 -175
rect 138 -177 140 -175
rect 143 -180 145 -175
rect 164 -180 166 -175
rect 180 -177 182 -175
rect 196 -177 198 -175
rect 201 -180 203 -175
rect 217 -177 219 -175
rect 233 -177 235 -175
rect 238 -178 240 -175
rect 254 -177 256 -175
rect 270 -177 272 -175
rect 275 -180 277 -175
rect 296 -180 298 -175
rect 312 -177 314 -175
rect 328 -177 330 -175
rect 333 -180 335 -175
rect 349 -177 351 -175
rect 365 -177 367 -175
rect 370 -178 372 -175
rect 386 -177 388 -175
rect 402 -177 404 -175
rect 407 -180 409 -175
rect 428 -180 430 -175
rect 444 -177 446 -175
rect 460 -177 462 -175
rect 465 -180 467 -175
rect 481 -177 483 -175
<< polycontact >>
rect 106 225 110 229
rect 143 225 147 229
rect 163 225 167 229
rect 201 225 205 229
rect 238 225 242 229
rect 275 225 279 229
rect 295 225 299 229
rect 333 225 337 229
rect 370 225 374 229
rect 407 225 411 229
rect 427 225 431 229
rect 465 225 469 229
rect 100 205 104 209
rect 118 207 122 211
rect 178 207 182 211
rect 136 198 140 205
rect 194 198 198 205
rect 213 202 217 206
rect 231 207 235 211
rect 250 207 254 211
rect 310 207 314 211
rect 268 198 272 205
rect 326 198 330 205
rect 345 202 349 206
rect 363 207 367 211
rect 382 207 386 211
rect 442 207 446 211
rect 400 198 404 205
rect 458 198 462 205
rect 479 202 483 206
rect 106 184 110 188
rect 143 182 147 186
rect 163 182 167 186
rect 199 182 203 186
rect 238 184 242 188
rect 275 182 279 186
rect 295 182 299 186
rect 331 182 335 186
rect 370 184 374 188
rect 407 182 411 186
rect 427 182 431 186
rect 463 182 467 186
rect 215 154 219 158
rect 239 154 243 158
rect 235 129 239 133
rect 250 121 254 125
rect 215 106 219 110
rect 239 106 243 110
rect 106 85 110 89
rect 143 85 147 89
rect 163 85 167 89
rect 201 85 205 89
rect 238 85 242 89
rect 275 85 279 89
rect 295 85 299 89
rect 333 85 337 89
rect 370 85 374 89
rect 407 85 411 89
rect 427 85 431 89
rect 465 85 469 89
rect 100 65 104 69
rect 118 67 122 71
rect 178 67 182 71
rect 136 58 140 65
rect 194 58 198 65
rect 213 62 217 66
rect 231 67 235 71
rect 250 67 254 71
rect 310 67 314 71
rect 268 58 272 65
rect 326 58 330 65
rect 345 62 349 66
rect 363 67 367 71
rect 382 67 386 71
rect 442 67 446 71
rect 400 58 404 65
rect 458 58 462 65
rect 479 62 483 66
rect 106 44 110 48
rect 143 42 147 46
rect 163 42 167 46
rect 199 42 203 46
rect 238 44 242 48
rect 275 42 279 46
rect 295 42 299 46
rect 331 42 335 46
rect 370 44 374 48
rect 407 42 411 46
rect 427 42 431 46
rect 463 42 467 46
rect 106 -1 110 3
rect 143 -1 147 3
rect 163 -1 167 3
rect 201 -1 205 3
rect 238 -1 242 3
rect 275 -1 279 3
rect 295 -1 299 3
rect 333 -1 337 3
rect 370 -1 374 3
rect 407 -1 411 3
rect 427 -1 431 3
rect 465 -1 469 3
rect 100 -21 104 -17
rect 118 -19 122 -15
rect 178 -19 182 -15
rect 136 -28 140 -21
rect 194 -28 198 -21
rect 213 -24 217 -20
rect 231 -19 235 -15
rect 250 -19 254 -15
rect 310 -19 314 -15
rect 268 -28 272 -21
rect 326 -28 330 -21
rect 345 -24 349 -20
rect 363 -19 367 -15
rect 382 -19 386 -15
rect 442 -19 446 -15
rect 400 -28 404 -21
rect 458 -28 462 -21
rect 479 -24 483 -20
rect 106 -42 110 -38
rect 143 -44 147 -40
rect 163 -44 167 -40
rect 199 -44 203 -40
rect 238 -42 242 -38
rect 275 -44 279 -40
rect 295 -44 299 -40
rect 331 -44 335 -40
rect 370 -42 374 -38
rect 407 -44 411 -40
rect 427 -44 431 -40
rect 463 -44 467 -40
rect 332 -72 336 -68
rect 356 -72 360 -68
rect 352 -97 356 -93
rect 367 -105 371 -101
rect 332 -120 336 -116
rect 356 -120 360 -116
rect 106 -141 110 -137
rect 143 -141 147 -137
rect 163 -141 167 -137
rect 201 -141 205 -137
rect 238 -141 242 -137
rect 275 -141 279 -137
rect 295 -141 299 -137
rect 333 -141 337 -137
rect 370 -141 374 -137
rect 407 -141 411 -137
rect 427 -141 431 -137
rect 465 -141 469 -137
rect 100 -161 104 -157
rect 118 -159 122 -155
rect 178 -159 182 -155
rect 136 -168 140 -161
rect 194 -168 198 -161
rect 213 -164 217 -160
rect 231 -159 235 -155
rect 250 -159 254 -155
rect 310 -159 314 -155
rect 268 -168 272 -161
rect 326 -168 330 -161
rect 345 -164 349 -160
rect 363 -159 367 -155
rect 382 -159 386 -155
rect 442 -159 446 -155
rect 400 -168 404 -161
rect 458 -168 462 -161
rect 479 -164 483 -160
rect 106 -182 110 -178
rect 143 -184 147 -180
rect 163 -184 167 -180
rect 199 -184 203 -180
rect 238 -182 242 -178
rect 275 -184 279 -180
rect 295 -184 299 -180
rect 331 -184 335 -180
rect 370 -182 374 -178
rect 407 -184 411 -180
rect 427 -184 431 -180
rect 463 -184 467 -180
<< metal1 >>
rect 93 239 102 243
rect 106 239 138 243
rect 142 239 205 243
rect 209 239 234 243
rect 238 239 270 243
rect 274 239 337 243
rect 341 239 366 243
rect 370 239 402 243
rect 406 239 469 243
rect 473 239 489 243
rect 93 232 126 236
rect 130 232 154 236
rect 158 232 184 236
rect 188 232 221 236
rect 225 232 258 236
rect 262 232 286 236
rect 290 232 316 236
rect 320 232 353 236
rect 357 232 390 236
rect 394 232 418 236
rect 422 232 448 236
rect 452 232 485 236
rect 96 222 99 232
rect 117 222 120 232
rect 133 222 136 232
rect 147 225 152 229
rect 156 225 163 229
rect 175 222 178 232
rect 191 222 194 232
rect 212 222 215 232
rect 228 222 231 232
rect 249 222 252 232
rect 265 222 268 232
rect 279 225 284 229
rect 288 225 295 229
rect 307 222 310 232
rect 323 222 326 232
rect 344 222 347 232
rect 360 222 363 232
rect 381 222 384 232
rect 397 222 400 232
rect 411 225 416 229
rect 420 225 427 229
rect 439 222 442 232
rect 455 222 458 232
rect 476 222 479 232
rect 113 208 118 211
rect 122 208 146 211
rect 171 208 178 211
rect 182 208 204 211
rect 224 208 231 211
rect 245 208 250 211
rect 254 208 278 211
rect 303 208 310 211
rect 314 208 336 211
rect 356 208 363 211
rect 377 208 382 211
rect 386 208 410 211
rect 435 208 442 211
rect 446 208 468 211
rect 129 198 136 201
rect 140 202 159 205
rect 159 195 162 201
rect 187 198 194 201
rect 198 202 213 205
rect 261 198 268 201
rect 272 202 291 205
rect 291 195 294 201
rect 319 198 326 201
rect 330 202 345 205
rect 393 198 400 201
rect 404 202 423 205
rect 423 195 426 201
rect 451 198 458 201
rect 462 202 479 205
rect 96 179 99 191
rect 117 179 120 191
rect 133 179 136 191
rect 147 182 159 185
rect 175 179 178 191
rect 191 179 194 191
rect 212 179 215 191
rect 228 179 231 191
rect 249 179 252 191
rect 265 179 268 191
rect 279 182 291 185
rect 307 179 310 191
rect 323 179 326 191
rect 344 179 347 191
rect 360 179 363 191
rect 381 179 384 191
rect 397 179 400 191
rect 411 182 423 185
rect 439 179 442 191
rect 455 179 458 191
rect 476 179 479 191
rect 93 175 126 179
rect 130 175 154 179
rect 158 175 184 179
rect 188 175 258 179
rect 262 175 286 179
rect 290 175 316 179
rect 320 175 390 179
rect 394 175 418 179
rect 422 175 448 179
rect 452 175 489 179
rect 93 168 102 172
rect 106 168 153 172
rect 157 168 203 172
rect 207 168 234 172
rect 238 168 285 172
rect 289 168 335 172
rect 339 168 366 172
rect 370 168 417 172
rect 421 168 467 172
rect 471 168 489 172
rect 100 162 484 165
rect 243 155 352 158
rect 223 147 227 151
rect 231 147 235 151
rect 79 136 211 140
rect 215 136 231 140
rect 247 136 502 140
rect 239 129 484 132
rect 254 122 484 125
rect 223 113 227 117
rect 231 113 235 117
rect 243 106 353 109
rect 93 99 102 103
rect 106 99 138 103
rect 142 99 205 103
rect 209 99 234 103
rect 238 99 270 103
rect 274 99 337 103
rect 341 99 366 103
rect 370 99 402 103
rect 406 99 469 103
rect 473 99 489 103
rect 93 92 126 96
rect 130 92 154 96
rect 158 92 184 96
rect 188 92 221 96
rect 225 92 258 96
rect 262 92 286 96
rect 290 92 316 96
rect 320 92 353 96
rect 357 92 390 96
rect 394 92 418 96
rect 422 92 448 96
rect 452 92 485 96
rect 96 82 99 92
rect 117 82 120 92
rect 133 82 136 92
rect 147 85 152 89
rect 156 85 163 89
rect 175 82 178 92
rect 191 82 194 92
rect 212 82 215 92
rect 228 82 231 92
rect 249 82 252 92
rect 265 82 268 92
rect 279 85 284 89
rect 288 85 295 89
rect 307 82 310 92
rect 323 82 326 92
rect 344 82 347 92
rect 360 82 363 92
rect 381 82 384 92
rect 397 82 400 92
rect 411 85 416 89
rect 420 85 427 89
rect 439 82 442 92
rect 455 82 458 92
rect 476 82 479 92
rect 113 68 118 71
rect 122 68 146 71
rect 171 68 178 71
rect 182 68 204 71
rect 224 68 231 71
rect 245 68 250 71
rect 254 68 278 71
rect 303 68 310 71
rect 314 68 336 71
rect 356 68 363 71
rect 377 68 382 71
rect 386 68 410 71
rect 435 68 442 71
rect 446 68 468 71
rect 129 58 136 61
rect 140 62 159 65
rect 159 55 162 61
rect 187 58 194 61
rect 198 62 213 65
rect 261 58 268 61
rect 272 62 291 65
rect 291 55 294 61
rect 319 58 326 61
rect 330 62 345 65
rect 393 58 400 61
rect 404 62 423 65
rect 423 55 426 61
rect 451 58 458 61
rect 462 62 479 65
rect 96 39 99 51
rect 117 39 120 51
rect 133 39 136 51
rect 147 42 159 45
rect 175 39 178 51
rect 191 39 194 51
rect 212 39 215 51
rect 228 39 231 51
rect 249 39 252 51
rect 265 39 268 51
rect 279 42 291 45
rect 307 39 310 51
rect 323 39 326 51
rect 344 39 347 51
rect 360 39 363 51
rect 381 39 384 51
rect 397 39 400 51
rect 411 42 423 45
rect 439 39 442 51
rect 455 39 458 51
rect 476 39 479 51
rect 93 35 126 39
rect 130 35 154 39
rect 158 35 184 39
rect 188 35 258 39
rect 262 35 286 39
rect 290 35 316 39
rect 320 35 390 39
rect 394 35 418 39
rect 422 35 448 39
rect 452 35 489 39
rect 93 28 102 32
rect 106 28 153 32
rect 157 28 203 32
rect 207 28 234 32
rect 238 28 285 32
rect 289 28 335 32
rect 339 28 366 32
rect 370 28 417 32
rect 421 28 467 32
rect 471 28 489 32
rect 99 21 484 24
rect 93 13 102 17
rect 106 13 138 17
rect 142 13 205 17
rect 209 13 234 17
rect 238 13 270 17
rect 274 13 337 17
rect 341 13 366 17
rect 370 13 402 17
rect 406 13 469 17
rect 473 13 489 17
rect 93 6 126 10
rect 130 6 154 10
rect 158 6 184 10
rect 188 6 221 10
rect 225 6 258 10
rect 262 6 286 10
rect 290 6 316 10
rect 320 6 353 10
rect 357 6 390 10
rect 394 6 418 10
rect 422 6 448 10
rect 452 6 485 10
rect 96 -4 99 6
rect 117 -4 120 6
rect 133 -4 136 6
rect 147 -1 152 3
rect 156 -1 163 3
rect 175 -4 178 6
rect 191 -4 194 6
rect 212 -4 215 6
rect 228 -4 231 6
rect 249 -4 252 6
rect 265 -4 268 6
rect 279 -1 284 3
rect 288 -1 295 3
rect 307 -4 310 6
rect 323 -4 326 6
rect 344 -4 347 6
rect 360 -4 363 6
rect 381 -4 384 6
rect 397 -4 400 6
rect 411 -1 416 3
rect 420 -1 427 3
rect 439 -4 442 6
rect 455 -4 458 6
rect 476 -4 479 6
rect 113 -18 118 -15
rect 122 -18 146 -15
rect 171 -18 178 -15
rect 182 -18 204 -15
rect 224 -18 231 -15
rect 245 -18 250 -15
rect 254 -18 278 -15
rect 303 -18 310 -15
rect 314 -18 336 -15
rect 356 -18 363 -15
rect 377 -18 382 -15
rect 386 -18 410 -15
rect 435 -18 442 -15
rect 446 -18 468 -15
rect 129 -28 136 -25
rect 140 -24 159 -21
rect 159 -31 162 -25
rect 187 -28 194 -25
rect 198 -24 213 -21
rect 261 -28 268 -25
rect 272 -24 291 -21
rect 291 -31 294 -25
rect 319 -28 326 -25
rect 330 -24 345 -21
rect 393 -28 400 -25
rect 404 -24 423 -21
rect 423 -31 426 -25
rect 451 -28 458 -25
rect 462 -24 479 -21
rect 96 -47 99 -35
rect 117 -47 120 -35
rect 133 -47 136 -35
rect 147 -44 159 -41
rect 175 -47 178 -35
rect 191 -47 194 -35
rect 212 -47 215 -35
rect 228 -47 231 -35
rect 249 -47 252 -35
rect 265 -47 268 -35
rect 279 -44 291 -41
rect 307 -47 310 -35
rect 323 -47 326 -35
rect 344 -47 347 -35
rect 360 -47 363 -35
rect 381 -47 384 -35
rect 397 -47 400 -35
rect 411 -44 423 -41
rect 439 -47 442 -35
rect 455 -47 458 -35
rect 476 -47 479 -35
rect 93 -51 126 -47
rect 130 -51 154 -47
rect 158 -51 184 -47
rect 188 -51 258 -47
rect 262 -51 286 -47
rect 290 -51 316 -47
rect 320 -51 390 -47
rect 394 -51 418 -47
rect 422 -51 448 -47
rect 452 -51 489 -47
rect 93 -58 102 -54
rect 106 -58 153 -54
rect 157 -58 203 -54
rect 207 -58 234 -54
rect 238 -58 285 -54
rect 289 -58 335 -54
rect 339 -58 366 -54
rect 370 -58 417 -54
rect 421 -58 467 -54
rect 471 -58 489 -54
rect 99 -64 484 -61
rect 224 -71 328 -68
rect 340 -79 344 -75
rect 348 -79 352 -75
rect 76 -90 328 -86
rect 332 -90 348 -86
rect 364 -90 510 -86
rect 356 -97 484 -94
rect 371 -104 484 -101
rect 340 -113 344 -109
rect 348 -113 352 -109
rect 224 -120 328 -117
rect 93 -127 102 -123
rect 106 -127 138 -123
rect 142 -127 205 -123
rect 209 -127 234 -123
rect 238 -127 270 -123
rect 274 -127 337 -123
rect 341 -127 366 -123
rect 370 -127 402 -123
rect 406 -127 469 -123
rect 473 -127 489 -123
rect 93 -134 126 -130
rect 130 -134 154 -130
rect 158 -134 184 -130
rect 188 -134 221 -130
rect 225 -134 258 -130
rect 262 -134 286 -130
rect 290 -134 316 -130
rect 320 -134 353 -130
rect 357 -134 390 -130
rect 394 -134 418 -130
rect 422 -134 448 -130
rect 452 -134 485 -130
rect 96 -144 99 -134
rect 117 -144 120 -134
rect 133 -144 136 -134
rect 147 -141 152 -137
rect 156 -141 163 -137
rect 175 -144 178 -134
rect 191 -144 194 -134
rect 212 -144 215 -134
rect 228 -144 231 -134
rect 249 -144 252 -134
rect 265 -144 268 -134
rect 279 -141 284 -137
rect 288 -141 295 -137
rect 307 -144 310 -134
rect 323 -144 326 -134
rect 344 -144 347 -134
rect 360 -144 363 -134
rect 381 -144 384 -134
rect 397 -144 400 -134
rect 411 -141 416 -137
rect 420 -141 427 -137
rect 439 -144 442 -134
rect 455 -144 458 -134
rect 476 -144 479 -134
rect 113 -158 118 -155
rect 122 -158 146 -155
rect 171 -158 178 -155
rect 182 -158 204 -155
rect 224 -158 231 -155
rect 245 -158 250 -155
rect 254 -158 278 -155
rect 303 -158 310 -155
rect 314 -158 336 -155
rect 356 -158 363 -155
rect 377 -158 382 -155
rect 386 -158 410 -155
rect 435 -158 442 -155
rect 446 -158 468 -155
rect 129 -168 136 -165
rect 140 -164 159 -161
rect 159 -171 162 -165
rect 187 -168 194 -165
rect 198 -164 213 -161
rect 261 -168 268 -165
rect 272 -164 291 -161
rect 291 -171 294 -165
rect 319 -168 326 -165
rect 330 -164 345 -161
rect 393 -168 400 -165
rect 404 -164 423 -161
rect 423 -171 426 -165
rect 451 -168 458 -165
rect 462 -164 479 -161
rect 96 -187 99 -175
rect 117 -187 120 -175
rect 133 -187 136 -175
rect 147 -184 159 -181
rect 175 -187 178 -175
rect 191 -187 194 -175
rect 212 -187 215 -175
rect 228 -187 231 -175
rect 249 -187 252 -175
rect 265 -187 268 -175
rect 279 -184 291 -181
rect 307 -187 310 -175
rect 323 -187 326 -175
rect 344 -187 347 -175
rect 360 -187 363 -175
rect 381 -187 384 -175
rect 397 -187 400 -175
rect 411 -184 423 -181
rect 439 -187 442 -175
rect 455 -187 458 -175
rect 476 -187 479 -175
rect 93 -191 126 -187
rect 130 -191 154 -187
rect 158 -191 184 -187
rect 188 -191 258 -187
rect 262 -191 286 -187
rect 290 -191 316 -187
rect 320 -191 390 -187
rect 394 -191 418 -187
rect 422 -191 448 -187
rect 452 -191 489 -187
rect 93 -198 102 -194
rect 106 -198 153 -194
rect 157 -198 203 -194
rect 207 -198 234 -194
rect 238 -198 285 -194
rect 289 -198 335 -194
rect 339 -198 366 -194
rect 370 -198 417 -194
rect 421 -198 467 -194
rect 471 -198 489 -194
<< m2contact >>
rect 102 239 106 243
rect 138 239 142 243
rect 205 239 209 243
rect 234 239 238 243
rect 270 239 274 243
rect 337 239 341 243
rect 366 239 370 243
rect 402 239 406 243
rect 469 239 473 243
rect 102 225 106 229
rect 152 225 156 229
rect 205 225 209 229
rect 234 225 238 229
rect 284 225 288 229
rect 337 225 341 229
rect 366 225 370 229
rect 416 225 420 229
rect 469 225 473 229
rect 125 214 129 218
rect 96 205 100 209
rect 109 208 113 214
rect 146 208 150 214
rect 159 210 163 214
rect 183 214 187 218
rect 257 214 261 218
rect 167 208 171 214
rect 204 208 208 214
rect 220 208 224 214
rect 241 208 245 214
rect 278 208 282 214
rect 291 210 295 214
rect 315 214 319 218
rect 389 214 393 218
rect 299 208 303 214
rect 336 208 340 214
rect 352 208 356 214
rect 373 208 377 214
rect 410 208 414 214
rect 423 210 427 214
rect 447 214 451 218
rect 431 208 435 214
rect 468 208 472 214
rect 484 210 488 214
rect 109 195 113 199
rect 125 195 129 201
rect 159 201 163 205
rect 146 195 150 199
rect 167 195 171 199
rect 183 195 187 201
rect 204 195 208 199
rect 220 195 224 199
rect 241 195 245 199
rect 257 195 261 201
rect 291 201 295 205
rect 278 195 282 199
rect 299 195 303 199
rect 315 195 319 201
rect 336 195 340 199
rect 352 195 356 199
rect 373 195 377 199
rect 389 195 393 201
rect 423 201 427 205
rect 410 195 414 199
rect 431 195 435 199
rect 447 195 451 201
rect 468 195 472 199
rect 484 195 488 199
rect 102 184 106 188
rect 139 182 143 186
rect 159 182 163 186
rect 203 182 207 186
rect 234 184 238 188
rect 271 182 275 186
rect 291 182 295 186
rect 335 182 339 186
rect 366 184 370 188
rect 403 182 407 186
rect 423 182 427 186
rect 467 182 471 186
rect 102 168 106 172
rect 153 168 157 172
rect 203 168 207 172
rect 234 168 238 172
rect 285 168 289 172
rect 335 168 339 172
rect 366 168 370 172
rect 417 168 421 172
rect 467 168 471 172
rect 96 161 100 165
rect 484 161 488 165
rect 219 154 224 158
rect 352 154 356 158
rect 227 147 231 151
rect 211 143 215 147
rect 243 143 247 147
rect 211 136 215 140
rect 243 136 247 140
rect 227 129 231 133
rect 484 129 488 133
rect 484 121 488 125
rect 211 117 215 121
rect 243 117 247 121
rect 227 113 231 117
rect 219 106 224 110
rect 353 106 357 110
rect 102 99 106 103
rect 138 99 142 103
rect 205 99 209 103
rect 234 99 238 103
rect 270 99 274 103
rect 337 99 341 103
rect 366 99 370 103
rect 402 99 406 103
rect 469 99 473 103
rect 102 85 106 89
rect 152 85 156 89
rect 205 85 209 89
rect 234 85 238 89
rect 284 85 288 89
rect 337 85 341 89
rect 366 85 370 89
rect 416 85 420 89
rect 469 85 473 89
rect 125 74 129 78
rect 96 65 100 69
rect 109 68 113 74
rect 146 68 150 74
rect 159 70 163 74
rect 183 74 187 78
rect 257 74 261 78
rect 167 68 171 74
rect 204 68 208 74
rect 220 68 224 74
rect 241 68 245 74
rect 278 68 282 74
rect 291 70 295 74
rect 315 74 319 78
rect 389 74 393 78
rect 299 68 303 74
rect 336 68 340 74
rect 352 68 356 74
rect 373 68 377 74
rect 410 68 414 74
rect 423 70 427 74
rect 447 74 451 78
rect 431 68 435 74
rect 468 68 472 74
rect 484 70 488 74
rect 109 55 113 59
rect 125 55 129 61
rect 159 61 163 65
rect 146 55 150 59
rect 167 55 171 59
rect 183 55 187 61
rect 204 55 208 59
rect 220 55 224 59
rect 241 55 245 59
rect 257 55 261 61
rect 291 61 295 65
rect 278 55 282 59
rect 299 55 303 59
rect 315 55 319 61
rect 336 55 340 59
rect 352 55 356 59
rect 373 55 377 59
rect 389 55 393 61
rect 423 61 427 65
rect 410 55 414 59
rect 431 55 435 59
rect 447 55 451 61
rect 468 55 472 59
rect 484 55 488 59
rect 102 44 106 48
rect 139 42 143 46
rect 159 42 163 46
rect 203 42 207 46
rect 234 44 238 48
rect 271 42 275 46
rect 291 42 295 46
rect 335 42 339 46
rect 366 44 370 48
rect 403 42 407 46
rect 423 42 427 46
rect 467 42 471 46
rect 102 28 106 32
rect 153 28 157 32
rect 203 28 207 32
rect 234 28 238 32
rect 285 28 289 32
rect 335 28 339 32
rect 366 28 370 32
rect 417 28 421 32
rect 467 28 471 32
rect 95 21 99 25
rect 484 21 488 25
rect 102 13 106 17
rect 138 13 142 17
rect 205 13 209 17
rect 234 13 238 17
rect 270 13 274 17
rect 337 13 341 17
rect 366 13 370 17
rect 402 13 406 17
rect 469 13 473 17
rect 102 -1 106 3
rect 152 -1 156 3
rect 205 -1 209 3
rect 234 -1 238 3
rect 284 -1 288 3
rect 337 -1 341 3
rect 366 -1 370 3
rect 416 -1 420 3
rect 469 -1 473 3
rect 125 -12 129 -8
rect 96 -21 100 -17
rect 109 -18 113 -12
rect 146 -18 150 -12
rect 159 -16 163 -12
rect 183 -12 187 -8
rect 257 -12 261 -8
rect 167 -18 171 -12
rect 204 -18 208 -12
rect 220 -18 224 -12
rect 241 -18 245 -12
rect 278 -18 282 -12
rect 291 -16 295 -12
rect 315 -12 319 -8
rect 389 -12 393 -8
rect 299 -18 303 -12
rect 336 -18 340 -12
rect 352 -18 356 -12
rect 373 -18 377 -12
rect 410 -18 414 -12
rect 423 -16 427 -12
rect 447 -12 451 -8
rect 431 -18 435 -12
rect 468 -18 472 -12
rect 484 -16 488 -12
rect 109 -31 113 -27
rect 125 -31 129 -25
rect 159 -25 163 -21
rect 146 -31 150 -27
rect 167 -31 171 -27
rect 183 -31 187 -25
rect 204 -31 208 -27
rect 220 -31 224 -27
rect 241 -31 245 -27
rect 257 -31 261 -25
rect 291 -25 295 -21
rect 278 -31 282 -27
rect 299 -31 303 -27
rect 315 -31 319 -25
rect 336 -31 340 -27
rect 352 -31 356 -27
rect 373 -31 377 -27
rect 389 -31 393 -25
rect 423 -25 427 -21
rect 410 -31 414 -27
rect 431 -31 435 -27
rect 447 -31 451 -25
rect 468 -31 472 -27
rect 484 -31 488 -27
rect 102 -42 106 -38
rect 139 -44 143 -40
rect 159 -44 163 -40
rect 203 -44 207 -40
rect 234 -42 238 -38
rect 271 -44 275 -40
rect 291 -44 295 -40
rect 335 -44 339 -40
rect 366 -42 370 -38
rect 403 -44 407 -40
rect 423 -44 427 -40
rect 467 -44 471 -40
rect 102 -58 106 -54
rect 153 -58 157 -54
rect 203 -58 207 -54
rect 234 -58 238 -54
rect 285 -58 289 -54
rect 335 -58 339 -54
rect 366 -58 370 -54
rect 417 -58 421 -54
rect 467 -58 471 -54
rect 95 -65 99 -61
rect 484 -65 488 -61
rect 220 -72 224 -68
rect 328 -72 332 -68
rect 352 -72 356 -68
rect 344 -79 348 -75
rect 328 -83 332 -79
rect 360 -83 364 -79
rect 328 -90 332 -86
rect 360 -90 364 -86
rect 344 -97 348 -93
rect 484 -97 488 -93
rect 484 -105 488 -101
rect 328 -109 332 -105
rect 360 -109 364 -105
rect 344 -113 348 -109
rect 220 -120 224 -116
rect 328 -120 332 -116
rect 352 -120 356 -116
rect 102 -127 106 -123
rect 138 -127 142 -123
rect 205 -127 209 -123
rect 234 -127 238 -123
rect 270 -127 274 -123
rect 337 -127 341 -123
rect 366 -127 370 -123
rect 402 -127 406 -123
rect 469 -127 473 -123
rect 102 -141 106 -137
rect 152 -141 156 -137
rect 205 -141 209 -137
rect 234 -141 238 -137
rect 284 -141 288 -137
rect 337 -141 341 -137
rect 366 -141 370 -137
rect 416 -141 420 -137
rect 469 -141 473 -137
rect 125 -152 129 -148
rect 96 -161 100 -157
rect 109 -158 113 -152
rect 146 -158 150 -152
rect 159 -156 163 -152
rect 183 -152 187 -148
rect 257 -152 261 -148
rect 167 -158 171 -152
rect 204 -158 208 -152
rect 220 -158 224 -152
rect 241 -158 245 -152
rect 278 -158 282 -152
rect 291 -156 295 -152
rect 315 -152 319 -148
rect 389 -152 393 -148
rect 299 -158 303 -152
rect 336 -158 340 -152
rect 352 -158 356 -152
rect 373 -158 377 -152
rect 410 -158 414 -152
rect 423 -156 427 -152
rect 447 -152 451 -148
rect 431 -158 435 -152
rect 468 -158 472 -152
rect 484 -156 488 -152
rect 109 -171 113 -167
rect 125 -171 129 -165
rect 159 -165 163 -161
rect 146 -171 150 -167
rect 167 -171 171 -167
rect 183 -171 187 -165
rect 204 -171 208 -167
rect 220 -171 224 -167
rect 241 -171 245 -167
rect 257 -171 261 -165
rect 291 -165 295 -161
rect 278 -171 282 -167
rect 299 -171 303 -167
rect 315 -171 319 -165
rect 336 -171 340 -167
rect 352 -171 356 -167
rect 373 -171 377 -167
rect 389 -171 393 -165
rect 423 -165 427 -161
rect 410 -171 414 -167
rect 431 -171 435 -167
rect 447 -171 451 -165
rect 468 -171 472 -167
rect 484 -171 488 -167
rect 102 -182 106 -178
rect 139 -184 143 -180
rect 159 -184 163 -180
rect 203 -184 207 -180
rect 234 -182 238 -178
rect 271 -184 275 -180
rect 291 -184 295 -180
rect 335 -184 339 -180
rect 366 -182 370 -178
rect 403 -184 407 -180
rect 423 -184 427 -180
rect 467 -184 471 -180
rect 102 -198 106 -194
rect 153 -198 157 -194
rect 203 -198 207 -194
rect 234 -198 238 -194
rect 285 -198 289 -194
rect 335 -198 339 -194
rect 366 -198 370 -194
rect 417 -198 421 -194
rect 467 -198 471 -194
<< metal2 >>
rect 103 229 106 239
rect 93 205 96 208
rect 110 199 113 208
rect 126 201 129 214
rect 139 186 142 239
rect 206 229 209 239
rect 146 214 150 218
rect 147 199 150 208
rect 102 172 105 184
rect 143 182 144 186
rect 153 172 156 225
rect 159 205 162 210
rect 168 199 171 208
rect 184 201 187 214
rect 205 199 208 208
rect 221 199 224 208
rect 204 172 207 182
rect 96 69 99 161
rect 221 158 224 195
rect 227 151 231 264
rect 235 229 238 239
rect 242 199 245 208
rect 258 201 261 214
rect 271 186 274 239
rect 338 229 341 239
rect 278 214 282 218
rect 279 199 282 208
rect 234 172 237 184
rect 275 182 276 186
rect 285 172 288 225
rect 291 205 294 210
rect 300 199 303 208
rect 316 201 319 214
rect 337 199 340 208
rect 336 172 339 182
rect 211 140 215 143
rect 211 121 215 136
rect 227 133 231 147
rect 243 147 247 151
rect 243 140 247 143
rect 243 121 247 136
rect 227 117 231 118
rect 243 113 247 117
rect 103 89 106 99
rect 110 59 113 68
rect 126 61 129 74
rect 139 46 142 99
rect 206 89 209 99
rect 146 74 150 78
rect 147 59 150 68
rect 102 32 105 44
rect 143 42 144 46
rect 153 32 156 85
rect 221 74 224 106
rect 159 65 162 70
rect 168 59 171 68
rect 184 61 187 74
rect 205 59 208 68
rect 221 59 224 68
rect 204 32 207 42
rect 96 -17 99 21
rect 103 3 106 13
rect 110 -27 113 -18
rect 126 -25 129 -12
rect 139 -40 142 13
rect 206 3 209 13
rect 146 -12 150 -8
rect 147 -27 150 -18
rect 102 -54 105 -42
rect 143 -44 144 -40
rect 153 -54 156 -1
rect 159 -21 162 -16
rect 168 -27 171 -18
rect 184 -25 187 -12
rect 205 -27 208 -18
rect 221 -27 224 -18
rect 204 -54 207 -44
rect 96 -157 99 -65
rect 221 -68 224 -31
rect 103 -137 106 -127
rect 110 -167 113 -158
rect 126 -165 129 -152
rect 139 -180 142 -127
rect 206 -137 209 -127
rect 146 -152 150 -148
rect 147 -167 150 -158
rect 102 -194 105 -182
rect 143 -184 144 -180
rect 153 -194 156 -141
rect 221 -152 224 -120
rect 159 -161 162 -156
rect 168 -167 171 -158
rect 184 -165 187 -152
rect 205 -167 208 -158
rect 221 -167 224 -158
rect 204 -194 207 -184
rect 227 -224 231 113
rect 235 89 238 99
rect 242 59 245 68
rect 258 61 261 74
rect 271 46 274 99
rect 338 89 341 99
rect 278 74 282 78
rect 279 59 282 68
rect 234 32 237 44
rect 275 42 276 46
rect 285 32 288 85
rect 291 65 294 70
rect 300 59 303 68
rect 316 61 319 74
rect 337 59 340 68
rect 336 32 339 42
rect 235 3 238 13
rect 242 -27 245 -18
rect 258 -25 261 -12
rect 271 -40 274 13
rect 338 3 341 13
rect 278 -12 282 -8
rect 279 -27 282 -18
rect 234 -54 237 -42
rect 275 -44 276 -40
rect 285 -54 288 -1
rect 291 -21 294 -16
rect 300 -27 303 -18
rect 316 -25 319 -12
rect 337 -27 340 -18
rect 336 -54 339 -44
rect 344 -75 348 261
rect 367 229 370 239
rect 353 199 356 208
rect 374 199 377 208
rect 390 201 393 214
rect 353 158 356 195
rect 403 186 406 239
rect 470 229 473 239
rect 410 214 414 218
rect 411 199 414 208
rect 366 172 369 184
rect 407 182 408 186
rect 417 172 420 225
rect 423 205 426 210
rect 432 199 435 208
rect 448 201 451 214
rect 469 199 472 208
rect 485 199 488 210
rect 468 172 471 182
rect 485 165 488 195
rect 485 133 488 161
rect 353 74 356 106
rect 367 89 370 99
rect 353 59 356 68
rect 374 59 377 68
rect 390 61 393 74
rect 403 46 406 99
rect 470 89 473 99
rect 410 74 414 78
rect 411 59 414 68
rect 366 32 369 44
rect 407 42 408 46
rect 417 32 420 85
rect 485 74 488 121
rect 423 65 426 70
rect 432 59 435 68
rect 448 61 451 74
rect 469 59 472 68
rect 485 59 488 70
rect 468 32 471 42
rect 485 25 488 55
rect 367 3 370 13
rect 353 -27 356 -18
rect 374 -27 377 -18
rect 390 -25 393 -12
rect 353 -68 356 -31
rect 403 -40 406 13
rect 470 3 473 13
rect 410 -12 414 -8
rect 411 -27 414 -18
rect 366 -54 369 -42
rect 407 -44 408 -40
rect 417 -54 420 -1
rect 423 -21 426 -16
rect 432 -27 435 -18
rect 448 -25 451 -12
rect 469 -27 472 -18
rect 485 -27 488 -16
rect 468 -54 471 -44
rect 485 -61 488 -31
rect 328 -86 332 -83
rect 328 -105 332 -90
rect 344 -93 348 -79
rect 360 -79 364 -75
rect 360 -86 364 -83
rect 360 -105 364 -90
rect 485 -93 488 -65
rect 344 -109 348 -108
rect 360 -113 364 -109
rect 235 -137 238 -127
rect 242 -167 245 -158
rect 258 -165 261 -152
rect 271 -180 274 -127
rect 338 -137 341 -127
rect 278 -152 282 -148
rect 279 -167 282 -158
rect 234 -194 237 -182
rect 275 -184 276 -180
rect 285 -194 288 -141
rect 291 -161 294 -156
rect 300 -167 303 -158
rect 316 -165 319 -152
rect 337 -167 340 -158
rect 336 -194 339 -184
rect 344 -222 348 -113
rect 353 -152 356 -120
rect 367 -137 370 -127
rect 353 -167 356 -158
rect 374 -167 377 -158
rect 390 -165 393 -152
rect 403 -180 406 -127
rect 470 -137 473 -127
rect 410 -152 414 -148
rect 411 -167 414 -158
rect 366 -194 369 -182
rect 407 -184 408 -180
rect 417 -194 420 -141
rect 485 -152 488 -105
rect 423 -161 426 -156
rect 432 -167 435 -158
rect 448 -165 451 -152
rect 469 -167 472 -158
rect 485 -167 488 -156
rect 468 -194 471 -184
<< labels >>
rlabel metal1 96 232 99 236 1 Vdd!
rlabel metal1 97 175 100 179 1 GND!
rlabel metal1 98 168 101 172 2 ~clk
rlabel metal1 96 239 99 243 4 clk
rlabel metal2 94 207 94 207 3 D
rlabel metal1 228 232 231 236 1 Vdd!
rlabel metal1 229 175 232 179 1 GND!
rlabel metal1 230 168 233 172 2 ~clk
rlabel metal1 228 239 231 243 4 clk
rlabel metal1 360 232 363 236 1 Vdd!
rlabel metal1 361 175 364 179 1 GND!
rlabel metal1 362 168 365 172 2 ~clk
rlabel metal1 360 239 363 243 4 clk
rlabel polysilicon 217 152 217 152 1 0
rlabel polysilicon 241 152 241 152 1 1
rlabel polysilicon 237 141 237 141 1 2
rlabel metal1 96 92 99 96 1 Vdd!
rlabel metal1 97 35 100 39 1 GND!
rlabel metal1 98 28 101 32 2 ~clk
rlabel metal1 96 99 99 103 4 clk
rlabel metal1 228 92 231 96 1 Vdd!
rlabel metal1 229 35 232 39 1 GND!
rlabel metal1 230 28 233 32 2 ~clk
rlabel metal1 228 99 231 103 4 clk
rlabel metal1 360 92 363 96 1 Vdd!
rlabel metal1 361 35 364 39 1 GND!
rlabel metal1 362 28 365 32 2 ~clk
rlabel metal1 360 99 363 103 4 clk
rlabel metal1 360 13 363 17 4 clk
rlabel metal1 362 -58 365 -54 2 ~clk
rlabel metal1 361 -51 364 -47 1 GND!
rlabel metal1 360 6 363 10 1 Vdd!
rlabel metal1 228 13 231 17 4 clk
rlabel metal1 230 -58 233 -54 2 ~clk
rlabel metal1 229 -51 232 -47 1 GND!
rlabel metal1 228 6 231 10 1 Vdd!
rlabel metal1 96 13 99 17 4 clk
rlabel metal1 98 -58 101 -54 2 ~clk
rlabel metal1 97 -51 100 -47 1 GND!
rlabel metal1 96 6 99 10 1 Vdd!
rlabel metal1 360 -127 363 -123 4 clk
rlabel metal1 362 -198 365 -194 2 ~clk
rlabel metal1 361 -191 364 -187 1 GND!
rlabel metal1 360 -134 363 -130 1 Vdd!
rlabel metal1 228 -127 231 -123 4 clk
rlabel metal1 230 -198 233 -194 2 ~clk
rlabel metal1 229 -191 232 -187 1 GND!
rlabel metal1 228 -134 231 -130 1 Vdd!
rlabel metal1 96 -127 99 -123 4 clk
rlabel metal1 98 -198 101 -194 2 ~clk
rlabel metal1 97 -191 100 -187 1 GND!
rlabel metal1 96 -134 99 -130 1 Vdd!
rlabel polysilicon 334 -73 334 -73 1 6
rlabel polysilicon 358 -73 358 -73 1 7
rlabel polysilicon 354 -91 354 -91 1 8
rlabel polysilicon 217 112 217 112 1 3
rlabel polysilicon 241 112 241 112 1 4
rlabel polysilicon 239 123 239 123 1 5
rlabel polysilicon 334 -114 334 -114 1 9
rlabel polysilicon 358 -115 358 -115 1 10
rlabel polysilicon 353 -103 353 -103 1 11
<< end >>
